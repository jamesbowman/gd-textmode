`default_nettype none

module top(
  input clka,
  output [2:0] vga_red,
  output [2:0] vga_green,
  output [2:0] vga_blue,
  output vga_hsync_n,
  output vga_vsync_n,

  input SCK,  // arduino 13
  input MOSI, // arduino 11
  output MISO, // arduino 12
  input SSEL, // arduino 9
  input AUX,  // arduino 2
  output AUDIOL,
  output AUDIOR,

  output flashMOSI,
  input  flashMISO,
  output flashSCK,
  output flashSSEL
  );

  wire ck_fb;
  wire clk;
  DCM #(
     .CLKFX_MULTIPLY(13),
     .CLKFX_DIVIDE(5),
     .DFS_FREQUENCY_MODE("LOW"), // HIGH or LOW frequency mode for frequency synthesis
     .DUTY_CYCLE_CORRECTION("TRUE"), // Duty cycle correction, TRUE or FALSE
     .STARTUP_WAIT("TRUE")    // Delay configuration DONE until DCM LOCK, TRUE/FALSE
  ) DCM_inst (
     .CLK0(ck_fb),    
     .CLKFX(clk), 
     .CLKFB(ck_fb),    // DCM clock feedback
     .CLKIN(clka),     // Clock input (from IBUFG, BUFG or DCM)
     .RST(0)
  );

  wire we;
  wire [7:0] wd;
  wire textMISO;

  spi _s (.clk(clk),
          .SCK(SCK),
          .MOSI(MOSI),
          .MISO(textMISO),
          .SSEL(SSEL),
          .we(we),
          .byte_recv(wd),
          .byte_xmit(8'ha0));

  reg[14:0] a;
  wire wclk = SCK;

  textmode tm(.wclk(wclk), 
              .write(we),
              .addr(a),
              .d(wd),
              .clk(clk),
              .vga_red(vga_red),
              .vga_green(vga_green),
              .vga_blue(vga_blue),
              .vga_hsync_n(vga_hsync_n),
              .vga_vsync_n(vga_vsync_n));

  always @(posedge SSEL or posedge SCK)
    if (SSEL == 1)
      a <= 5;
    else if (we)
      a <= a + 1;

  assign AUDIOL = 0;
  assign AUDIOR = 0;

  assign flashMOSI = MOSI;
  assign flashSCK = SCK;
  assign flashSSEL = AUX;

  assign MISO = (SSEL == 0) ? textMISO : flashMISO;

endmodule

module spi(
  input clk,
  input SCK, input MOSI, output MISO, input SSEL,

  output we,
  output [7:0] byte_recv,
  input [7:0] byte_xmit);

  reg [2:0] bit;
  reg [7:0] recv;
  wire [7:0] recvN = {recv[6:0], MOSI};

  always @(posedge SSEL or posedge SCK)
    if (SSEL == 1)
      bit <= 7;
    else begin
      recv <= recvN;
      bit <= bit - 1;
    end

  assign MISO = byte_xmit[bit[2:0]];
  assign byte_recv = recvN;
  assign we = !SSEL & (bit == 0);
endmodule

module ram16k(
    input           wclk,
    input           We,
    input  [13:0]    Waddr,
    input  [7:0]   Din,

    input           rclk,
    input  [13:0]    Raddr,
    output [7:0]   Dout);
 
    //synthesis attribute ram_style of mem is block
    reg    [7:0]  mem[0:16383]; //pragma attribute mem ram_block TRUE
    reg    [13:0]  raddr_reg;
 
    initial begin
        $readmemh("init.hex", mem);
    end

    always @ (posedge wclk)
      if (We)
        mem[Waddr]  <= Din;  
 
    always @ (posedge rclk)
      raddr_reg  <= Raddr;
      // Dout  <= mem[raddr_reg];   //registered read
 
    assign Dout = mem[raddr_reg];  //unregistered read            

endmodule

module textmode(
  input wclk,
  input write,
  input [14:0] addr,
  input [7:0] d,

  input clk,
  output reg [2:0] vga_red,
  output reg [2:0] vga_green,
  output reg [2:0] vga_blue,
  output reg vga_hsync_n,
  output reg vga_vsync_n);

  // http://tinyvga.com/vga-timing/1024x768@60Hz

  // hcounter:
  //  0   -1023   visible area
  //  1024-1047   front porch
  //  1048-1183   sync pulse
  //  1184-1343   back porch

  reg [10:0] hcounter;
  wire [10:0] hcounterN = (hcounter == 11'd1343) ? 11'd0 : (hcounter + 11'd1);

  // vcounter:
  //  0  -767     visble area
  //  768-770     front porch
  //  771-776     sync pulse
  //  777-805     back porch

  reg [9:0] vcounter;
  reg [9:0] vcounterN;
  always @*
    if (hcounterN != 11'd0)
      vcounterN = vcounter;
    else if (vcounter != 10'd805)
      vcounterN = vcounter + 1;
    else
      vcounterN = 10'd0;

  wire visible = (hcounter < 1024) & (vcounter < 768);

  wire [7:0] cc;
  ram16k r(.wclk(wclk), .rclk(clk), .We(write), .Waddr(addr[13:0]), .Raddr(hcounterN[10:3]), .Din(d), .Dout(cc));
  // assign cc = hcounterN[10:3] + vcounterN[9:4];
  wire pix;
  fontrom fr(.clk(clk), .ch(cc), .row(vcounterN[3:0]), .col(hcounterN[2:0] - 1), .pix(pix));

  always @(posedge clk) begin
    hcounter <= hcounterN;
    vcounter <= vcounterN;
    vga_hsync_n <= !((1048 <= hcounter) & (hcounter < 1184));
    vga_vsync_n <= !((771 <= vcounter) & (vcounter < 777));
    vga_red <= visible ? {pix, pix, pix} : 3'b000;
    vga_green <= visible ? {pix, pix, pix} : 3'b000;
    vga_blue <= visible ? {pix, pix, pix} : 3'b000;
  end
endmodule

module fontrom(
  input clk,
  input [7:0] ch,
  input [3:0] row,
  input [2:0] col,
  output pix);

  reg [11:0] a;
  reg [2:0] col_;
  always @(posedge clk) begin
    a <= {ch, row};
    col_ <= col;
  end
    
  reg [7:0] pattern;
  assign pix = pattern[~col_];
  always @*
  case (a)
    { 8'h00, 4'h0 }: pattern = 8'b00000000; 
    { 8'h00, 4'h1 }: pattern = 8'b00000000; 
    { 8'h00, 4'h2 }: pattern = 8'b00000000; 
    { 8'h00, 4'h3 }: pattern = 8'b00000000; 
    { 8'h00, 4'h4 }: pattern = 8'b00000000; 
    { 8'h00, 4'h5 }: pattern = 8'b00000000; 
    { 8'h00, 4'h6 }: pattern = 8'b00000000; 
    { 8'h00, 4'h7 }: pattern = 8'b00000000; 
    { 8'h00, 4'h8 }: pattern = 8'b00000000; 
    { 8'h00, 4'h9 }: pattern = 8'b00000000; 
    { 8'h00, 4'ha }: pattern = 8'b00000000; 
    { 8'h00, 4'hb }: pattern = 8'b00000000; 
    { 8'h00, 4'hc }: pattern = 8'b00000000; 
    { 8'h00, 4'hd }: pattern = 8'b00000000; 
    { 8'h00, 4'he }: pattern = 8'b00000000; 
    { 8'h00, 4'hf }: pattern = 8'b00000000; 

    { 8'h01, 4'h0 }: pattern = 8'b00000000; 
    { 8'h01, 4'h1 }: pattern = 8'b00000000; 
    { 8'h01, 4'h2 }: pattern = 8'b01111110; 
    { 8'h01, 4'h3 }: pattern = 8'b10000001; 
    { 8'h01, 4'h4 }: pattern = 8'b10100101; 
    { 8'h01, 4'h5 }: pattern = 8'b10000001; 
    { 8'h01, 4'h6 }: pattern = 8'b10000001; 
    { 8'h01, 4'h7 }: pattern = 8'b10111101; 
    { 8'h01, 4'h8 }: pattern = 8'b10011001; 
    { 8'h01, 4'h9 }: pattern = 8'b10000001; 
    { 8'h01, 4'ha }: pattern = 8'b10000001; 
    { 8'h01, 4'hb }: pattern = 8'b01111110; 
    { 8'h01, 4'hc }: pattern = 8'b00000000; 
    { 8'h01, 4'hd }: pattern = 8'b00000000; 
    { 8'h01, 4'he }: pattern = 8'b00000000; 
    { 8'h01, 4'hf }: pattern = 8'b00000000; 

    { 8'h02, 4'h0 }: pattern = 8'b00000000; 
    { 8'h02, 4'h1 }: pattern = 8'b00000000; 
    { 8'h02, 4'h2 }: pattern = 8'b01111110; 
    { 8'h02, 4'h3 }: pattern = 8'b11111111; 
    { 8'h02, 4'h4 }: pattern = 8'b11011011; 
    { 8'h02, 4'h5 }: pattern = 8'b11111111; 
    { 8'h02, 4'h6 }: pattern = 8'b11111111; 
    { 8'h02, 4'h7 }: pattern = 8'b11000011; 
    { 8'h02, 4'h8 }: pattern = 8'b11100111; 
    { 8'h02, 4'h9 }: pattern = 8'b11111111; 
    { 8'h02, 4'ha }: pattern = 8'b11111111; 
    { 8'h02, 4'hb }: pattern = 8'b01111110; 
    { 8'h02, 4'hc }: pattern = 8'b00000000; 
    { 8'h02, 4'hd }: pattern = 8'b00000000; 
    { 8'h02, 4'he }: pattern = 8'b00000000; 
    { 8'h02, 4'hf }: pattern = 8'b00000000; 

    { 8'h03, 4'h0 }: pattern = 8'b00000000; 
    { 8'h03, 4'h1 }: pattern = 8'b00000000; 
    { 8'h03, 4'h2 }: pattern = 8'b00000000; 
    { 8'h03, 4'h3 }: pattern = 8'b00000000; 
    { 8'h03, 4'h4 }: pattern = 8'b01101100; 
    { 8'h03, 4'h5 }: pattern = 8'b11111110; 
    { 8'h03, 4'h6 }: pattern = 8'b11111110; 
    { 8'h03, 4'h7 }: pattern = 8'b11111110; 
    { 8'h03, 4'h8 }: pattern = 8'b11111110; 
    { 8'h03, 4'h9 }: pattern = 8'b01111100; 
    { 8'h03, 4'ha }: pattern = 8'b00111000; 
    { 8'h03, 4'hb }: pattern = 8'b00010000; 
    { 8'h03, 4'hc }: pattern = 8'b00000000; 
    { 8'h03, 4'hd }: pattern = 8'b00000000; 
    { 8'h03, 4'he }: pattern = 8'b00000000; 
    { 8'h03, 4'hf }: pattern = 8'b00000000; 

    { 8'h04, 4'h0 }: pattern = 8'b00000000; 
    { 8'h04, 4'h1 }: pattern = 8'b00000000; 
    { 8'h04, 4'h2 }: pattern = 8'b00000000; 
    { 8'h04, 4'h3 }: pattern = 8'b00000000; 
    { 8'h04, 4'h4 }: pattern = 8'b00010000; 
    { 8'h04, 4'h5 }: pattern = 8'b00111000; 
    { 8'h04, 4'h6 }: pattern = 8'b01111100; 
    { 8'h04, 4'h7 }: pattern = 8'b11111110; 
    { 8'h04, 4'h8 }: pattern = 8'b01111100; 
    { 8'h04, 4'h9 }: pattern = 8'b00111000; 
    { 8'h04, 4'ha }: pattern = 8'b00010000; 
    { 8'h04, 4'hb }: pattern = 8'b00000000; 
    { 8'h04, 4'hc }: pattern = 8'b00000000; 
    { 8'h04, 4'hd }: pattern = 8'b00000000; 
    { 8'h04, 4'he }: pattern = 8'b00000000; 
    { 8'h04, 4'hf }: pattern = 8'b00000000; 

    { 8'h05, 4'h0 }: pattern = 8'b00000000; 
    { 8'h05, 4'h1 }: pattern = 8'b00000000; 
    { 8'h05, 4'h2 }: pattern = 8'b00000000; 
    { 8'h05, 4'h3 }: pattern = 8'b00011000; 
    { 8'h05, 4'h4 }: pattern = 8'b00111100; 
    { 8'h05, 4'h5 }: pattern = 8'b00111100; 
    { 8'h05, 4'h6 }: pattern = 8'b11100111; 
    { 8'h05, 4'h7 }: pattern = 8'b11100111; 
    { 8'h05, 4'h8 }: pattern = 8'b11100111; 
    { 8'h05, 4'h9 }: pattern = 8'b00011000; 
    { 8'h05, 4'ha }: pattern = 8'b00011000; 
    { 8'h05, 4'hb }: pattern = 8'b00111100; 
    { 8'h05, 4'hc }: pattern = 8'b00000000; 
    { 8'h05, 4'hd }: pattern = 8'b00000000; 
    { 8'h05, 4'he }: pattern = 8'b00000000; 
    { 8'h05, 4'hf }: pattern = 8'b00000000; 

    { 8'h06, 4'h0 }: pattern = 8'b00000000; 
    { 8'h06, 4'h1 }: pattern = 8'b00000000; 
    { 8'h06, 4'h2 }: pattern = 8'b00000000; 
    { 8'h06, 4'h3 }: pattern = 8'b00011000; 
    { 8'h06, 4'h4 }: pattern = 8'b00111100; 
    { 8'h06, 4'h5 }: pattern = 8'b01111110; 
    { 8'h06, 4'h6 }: pattern = 8'b11111111; 
    { 8'h06, 4'h7 }: pattern = 8'b11111111; 
    { 8'h06, 4'h8 }: pattern = 8'b01111110; 
    { 8'h06, 4'h9 }: pattern = 8'b00011000; 
    { 8'h06, 4'ha }: pattern = 8'b00011000; 
    { 8'h06, 4'hb }: pattern = 8'b00111100; 
    { 8'h06, 4'hc }: pattern = 8'b00000000; 
    { 8'h06, 4'hd }: pattern = 8'b00000000; 
    { 8'h06, 4'he }: pattern = 8'b00000000; 
    { 8'h06, 4'hf }: pattern = 8'b00000000; 

    { 8'h07, 4'h0 }: pattern = 8'b00000000; 
    { 8'h07, 4'h1 }: pattern = 8'b00000000; 
    { 8'h07, 4'h2 }: pattern = 8'b00000000; 
    { 8'h07, 4'h3 }: pattern = 8'b00000000; 
    { 8'h07, 4'h4 }: pattern = 8'b00000000; 
    { 8'h07, 4'h5 }: pattern = 8'b00000000; 
    { 8'h07, 4'h6 }: pattern = 8'b00011000; 
    { 8'h07, 4'h7 }: pattern = 8'b00111100; 
    { 8'h07, 4'h8 }: pattern = 8'b00111100; 
    { 8'h07, 4'h9 }: pattern = 8'b00011000; 
    { 8'h07, 4'ha }: pattern = 8'b00000000; 
    { 8'h07, 4'hb }: pattern = 8'b00000000; 
    { 8'h07, 4'hc }: pattern = 8'b00000000; 
    { 8'h07, 4'hd }: pattern = 8'b00000000; 
    { 8'h07, 4'he }: pattern = 8'b00000000; 
    { 8'h07, 4'hf }: pattern = 8'b00000000; 

    { 8'h08, 4'h0 }: pattern = 8'b11111111; 
    { 8'h08, 4'h1 }: pattern = 8'b11111111; 
    { 8'h08, 4'h2 }: pattern = 8'b11111111; 
    { 8'h08, 4'h3 }: pattern = 8'b11111111; 
    { 8'h08, 4'h4 }: pattern = 8'b11111111; 
    { 8'h08, 4'h5 }: pattern = 8'b11111111; 
    { 8'h08, 4'h6 }: pattern = 8'b11100111; 
    { 8'h08, 4'h7 }: pattern = 8'b11000011; 
    { 8'h08, 4'h8 }: pattern = 8'b11000011; 
    { 8'h08, 4'h9 }: pattern = 8'b11100111; 
    { 8'h08, 4'ha }: pattern = 8'b11111111; 
    { 8'h08, 4'hb }: pattern = 8'b11111111; 
    { 8'h08, 4'hc }: pattern = 8'b11111111; 
    { 8'h08, 4'hd }: pattern = 8'b11111111; 
    { 8'h08, 4'he }: pattern = 8'b11111111; 
    { 8'h08, 4'hf }: pattern = 8'b11111111; 

    { 8'h09, 4'h0 }: pattern = 8'b00000000; 
    { 8'h09, 4'h1 }: pattern = 8'b00000000; 
    { 8'h09, 4'h2 }: pattern = 8'b00000000; 
    { 8'h09, 4'h3 }: pattern = 8'b00000000; 
    { 8'h09, 4'h4 }: pattern = 8'b00000000; 
    { 8'h09, 4'h5 }: pattern = 8'b00111100; 
    { 8'h09, 4'h6 }: pattern = 8'b01100110; 
    { 8'h09, 4'h7 }: pattern = 8'b01000010; 
    { 8'h09, 4'h8 }: pattern = 8'b01000010; 
    { 8'h09, 4'h9 }: pattern = 8'b01100110; 
    { 8'h09, 4'ha }: pattern = 8'b00111100; 
    { 8'h09, 4'hb }: pattern = 8'b00000000; 
    { 8'h09, 4'hc }: pattern = 8'b00000000; 
    { 8'h09, 4'hd }: pattern = 8'b00000000; 
    { 8'h09, 4'he }: pattern = 8'b00000000; 
    { 8'h09, 4'hf }: pattern = 8'b00000000; 

    { 8'h0a, 4'h0 }: pattern = 8'b11111111; 
    { 8'h0a, 4'h1 }: pattern = 8'b11111111; 
    { 8'h0a, 4'h2 }: pattern = 8'b11111111; 
    { 8'h0a, 4'h3 }: pattern = 8'b11111111; 
    { 8'h0a, 4'h4 }: pattern = 8'b11111111; 
    { 8'h0a, 4'h5 }: pattern = 8'b11000011; 
    { 8'h0a, 4'h6 }: pattern = 8'b10011001; 
    { 8'h0a, 4'h7 }: pattern = 8'b10111101; 
    { 8'h0a, 4'h8 }: pattern = 8'b10111101; 
    { 8'h0a, 4'h9 }: pattern = 8'b10011001; 
    { 8'h0a, 4'ha }: pattern = 8'b11000011; 
    { 8'h0a, 4'hb }: pattern = 8'b11111111; 
    { 8'h0a, 4'hc }: pattern = 8'b11111111; 
    { 8'h0a, 4'hd }: pattern = 8'b11111111; 
    { 8'h0a, 4'he }: pattern = 8'b11111111; 
    { 8'h0a, 4'hf }: pattern = 8'b11111111; 

    { 8'h0b, 4'h0 }: pattern = 8'b00000000; 
    { 8'h0b, 4'h1 }: pattern = 8'b00000000; 
    { 8'h0b, 4'h2 }: pattern = 8'b00011110; 
    { 8'h0b, 4'h3 }: pattern = 8'b00001110; 
    { 8'h0b, 4'h4 }: pattern = 8'b00011010; 
    { 8'h0b, 4'h5 }: pattern = 8'b00110010; 
    { 8'h0b, 4'h6 }: pattern = 8'b01111000; 
    { 8'h0b, 4'h7 }: pattern = 8'b11001100; 
    { 8'h0b, 4'h8 }: pattern = 8'b11001100; 
    { 8'h0b, 4'h9 }: pattern = 8'b11001100; 
    { 8'h0b, 4'ha }: pattern = 8'b11001100; 
    { 8'h0b, 4'hb }: pattern = 8'b01111000; 
    { 8'h0b, 4'hc }: pattern = 8'b00000000; 
    { 8'h0b, 4'hd }: pattern = 8'b00000000; 
    { 8'h0b, 4'he }: pattern = 8'b00000000; 
    { 8'h0b, 4'hf }: pattern = 8'b00000000; 

    { 8'h0c, 4'h0 }: pattern = 8'b00000000; 
    { 8'h0c, 4'h1 }: pattern = 8'b00000000; 
    { 8'h0c, 4'h2 }: pattern = 8'b00111100; 
    { 8'h0c, 4'h3 }: pattern = 8'b01100110; 
    { 8'h0c, 4'h4 }: pattern = 8'b01100110; 
    { 8'h0c, 4'h5 }: pattern = 8'b01100110; 
    { 8'h0c, 4'h6 }: pattern = 8'b01100110; 
    { 8'h0c, 4'h7 }: pattern = 8'b00111100; 
    { 8'h0c, 4'h8 }: pattern = 8'b00011000; 
    { 8'h0c, 4'h9 }: pattern = 8'b01111110; 
    { 8'h0c, 4'ha }: pattern = 8'b00011000; 
    { 8'h0c, 4'hb }: pattern = 8'b00011000; 
    { 8'h0c, 4'hc }: pattern = 8'b00000000; 
    { 8'h0c, 4'hd }: pattern = 8'b00000000; 
    { 8'h0c, 4'he }: pattern = 8'b00000000; 
    { 8'h0c, 4'hf }: pattern = 8'b00000000; 

    { 8'h0d, 4'h0 }: pattern = 8'b00000000; 
    { 8'h0d, 4'h1 }: pattern = 8'b00000000; 
    { 8'h0d, 4'h2 }: pattern = 8'b00111111; 
    { 8'h0d, 4'h3 }: pattern = 8'b00110011; 
    { 8'h0d, 4'h4 }: pattern = 8'b00111111; 
    { 8'h0d, 4'h5 }: pattern = 8'b00110000; 
    { 8'h0d, 4'h6 }: pattern = 8'b00110000; 
    { 8'h0d, 4'h7 }: pattern = 8'b00110000; 
    { 8'h0d, 4'h8 }: pattern = 8'b00110000; 
    { 8'h0d, 4'h9 }: pattern = 8'b01110000; 
    { 8'h0d, 4'ha }: pattern = 8'b11110000; 
    { 8'h0d, 4'hb }: pattern = 8'b11100000; 
    { 8'h0d, 4'hc }: pattern = 8'b00000000; 
    { 8'h0d, 4'hd }: pattern = 8'b00000000; 
    { 8'h0d, 4'he }: pattern = 8'b00000000; 
    { 8'h0d, 4'hf }: pattern = 8'b00000000; 

    { 8'h0e, 4'h0 }: pattern = 8'b00000000; 
    { 8'h0e, 4'h1 }: pattern = 8'b00000000; 
    { 8'h0e, 4'h2 }: pattern = 8'b01111111; 
    { 8'h0e, 4'h3 }: pattern = 8'b01100011; 
    { 8'h0e, 4'h4 }: pattern = 8'b01111111; 
    { 8'h0e, 4'h5 }: pattern = 8'b01100011; 
    { 8'h0e, 4'h6 }: pattern = 8'b01100011; 
    { 8'h0e, 4'h7 }: pattern = 8'b01100011; 
    { 8'h0e, 4'h8 }: pattern = 8'b01100011; 
    { 8'h0e, 4'h9 }: pattern = 8'b01100111; 
    { 8'h0e, 4'ha }: pattern = 8'b11100111; 
    { 8'h0e, 4'hb }: pattern = 8'b11100110; 
    { 8'h0e, 4'hc }: pattern = 8'b11000000; 
    { 8'h0e, 4'hd }: pattern = 8'b00000000; 
    { 8'h0e, 4'he }: pattern = 8'b00000000; 
    { 8'h0e, 4'hf }: pattern = 8'b00000000; 

    { 8'h0f, 4'h0 }: pattern = 8'b00000000; 
    { 8'h0f, 4'h1 }: pattern = 8'b00000000; 
    { 8'h0f, 4'h2 }: pattern = 8'b00000000; 
    { 8'h0f, 4'h3 }: pattern = 8'b00011000; 
    { 8'h0f, 4'h4 }: pattern = 8'b00011000; 
    { 8'h0f, 4'h5 }: pattern = 8'b11011011; 
    { 8'h0f, 4'h6 }: pattern = 8'b00111100; 
    { 8'h0f, 4'h7 }: pattern = 8'b11100111; 
    { 8'h0f, 4'h8 }: pattern = 8'b00111100; 
    { 8'h0f, 4'h9 }: pattern = 8'b11011011; 
    { 8'h0f, 4'ha }: pattern = 8'b00011000; 
    { 8'h0f, 4'hb }: pattern = 8'b00011000; 
    { 8'h0f, 4'hc }: pattern = 8'b00000000; 
    { 8'h0f, 4'hd }: pattern = 8'b00000000; 
    { 8'h0f, 4'he }: pattern = 8'b00000000; 
    { 8'h0f, 4'hf }: pattern = 8'b00000000; 

    { 8'h10, 4'h0 }: pattern = 8'b00000000; 
    { 8'h10, 4'h1 }: pattern = 8'b10000000; 
    { 8'h10, 4'h2 }: pattern = 8'b11000000; 
    { 8'h10, 4'h3 }: pattern = 8'b11100000; 
    { 8'h10, 4'h4 }: pattern = 8'b11110000; 
    { 8'h10, 4'h5 }: pattern = 8'b11111000; 
    { 8'h10, 4'h6 }: pattern = 8'b11111110; 
    { 8'h10, 4'h7 }: pattern = 8'b11111000; 
    { 8'h10, 4'h8 }: pattern = 8'b11110000; 
    { 8'h10, 4'h9 }: pattern = 8'b11100000; 
    { 8'h10, 4'ha }: pattern = 8'b11000000; 
    { 8'h10, 4'hb }: pattern = 8'b10000000; 
    { 8'h10, 4'hc }: pattern = 8'b00000000; 
    { 8'h10, 4'hd }: pattern = 8'b00000000; 
    { 8'h10, 4'he }: pattern = 8'b00000000; 
    { 8'h10, 4'hf }: pattern = 8'b00000000; 

    { 8'h11, 4'h0 }: pattern = 8'b00000000; 
    { 8'h11, 4'h1 }: pattern = 8'b00000010; 
    { 8'h11, 4'h2 }: pattern = 8'b00000110; 
    { 8'h11, 4'h3 }: pattern = 8'b00001110; 
    { 8'h11, 4'h4 }: pattern = 8'b00011110; 
    { 8'h11, 4'h5 }: pattern = 8'b00111110; 
    { 8'h11, 4'h6 }: pattern = 8'b11111110; 
    { 8'h11, 4'h7 }: pattern = 8'b00111110; 
    { 8'h11, 4'h8 }: pattern = 8'b00011110; 
    { 8'h11, 4'h9 }: pattern = 8'b00001110; 
    { 8'h11, 4'ha }: pattern = 8'b00000110; 
    { 8'h11, 4'hb }: pattern = 8'b00000010; 
    { 8'h11, 4'hc }: pattern = 8'b00000000; 
    { 8'h11, 4'hd }: pattern = 8'b00000000; 
    { 8'h11, 4'he }: pattern = 8'b00000000; 
    { 8'h11, 4'hf }: pattern = 8'b00000000; 

    { 8'h12, 4'h0 }: pattern = 8'b00000000; 
    { 8'h12, 4'h1 }: pattern = 8'b00000000; 
    { 8'h12, 4'h2 }: pattern = 8'b00011000; 
    { 8'h12, 4'h3 }: pattern = 8'b00111100; 
    { 8'h12, 4'h4 }: pattern = 8'b01111110; 
    { 8'h12, 4'h5 }: pattern = 8'b00011000; 
    { 8'h12, 4'h6 }: pattern = 8'b00011000; 
    { 8'h12, 4'h7 }: pattern = 8'b00011000; 
    { 8'h12, 4'h8 }: pattern = 8'b01111110; 
    { 8'h12, 4'h9 }: pattern = 8'b00111100; 
    { 8'h12, 4'ha }: pattern = 8'b00011000; 
    { 8'h12, 4'hb }: pattern = 8'b00000000; 
    { 8'h12, 4'hc }: pattern = 8'b00000000; 
    { 8'h12, 4'hd }: pattern = 8'b00000000; 
    { 8'h12, 4'he }: pattern = 8'b00000000; 
    { 8'h12, 4'hf }: pattern = 8'b00000000; 

    { 8'h13, 4'h0 }: pattern = 8'b00000000; 
    { 8'h13, 4'h1 }: pattern = 8'b00000000; 
    { 8'h13, 4'h2 }: pattern = 8'b01100110; 
    { 8'h13, 4'h3 }: pattern = 8'b01100110; 
    { 8'h13, 4'h4 }: pattern = 8'b01100110; 
    { 8'h13, 4'h5 }: pattern = 8'b01100110; 
    { 8'h13, 4'h6 }: pattern = 8'b01100110; 
    { 8'h13, 4'h7 }: pattern = 8'b01100110; 
    { 8'h13, 4'h8 }: pattern = 8'b01100110; 
    { 8'h13, 4'h9 }: pattern = 8'b00000000; 
    { 8'h13, 4'ha }: pattern = 8'b01100110; 
    { 8'h13, 4'hb }: pattern = 8'b01100110; 
    { 8'h13, 4'hc }: pattern = 8'b00000000; 
    { 8'h13, 4'hd }: pattern = 8'b00000000; 
    { 8'h13, 4'he }: pattern = 8'b00000000; 
    { 8'h13, 4'hf }: pattern = 8'b00000000; 

    { 8'h14, 4'h0 }: pattern = 8'b00000000; 
    { 8'h14, 4'h1 }: pattern = 8'b00000000; 
    { 8'h14, 4'h2 }: pattern = 8'b01111111; 
    { 8'h14, 4'h3 }: pattern = 8'b11011011; 
    { 8'h14, 4'h4 }: pattern = 8'b11011011; 
    { 8'h14, 4'h5 }: pattern = 8'b11011011; 
    { 8'h14, 4'h6 }: pattern = 8'b01111011; 
    { 8'h14, 4'h7 }: pattern = 8'b00011011; 
    { 8'h14, 4'h8 }: pattern = 8'b00011011; 
    { 8'h14, 4'h9 }: pattern = 8'b00011011; 
    { 8'h14, 4'ha }: pattern = 8'b00011011; 
    { 8'h14, 4'hb }: pattern = 8'b00011011; 
    { 8'h14, 4'hc }: pattern = 8'b00000000; 
    { 8'h14, 4'hd }: pattern = 8'b00000000; 
    { 8'h14, 4'he }: pattern = 8'b00000000; 
    { 8'h14, 4'hf }: pattern = 8'b00000000; 

    { 8'h15, 4'h0 }: pattern = 8'b00000000; 
    { 8'h15, 4'h1 }: pattern = 8'b01111100; 
    { 8'h15, 4'h2 }: pattern = 8'b11000110; 
    { 8'h15, 4'h3 }: pattern = 8'b01100000; 
    { 8'h15, 4'h4 }: pattern = 8'b00111000; 
    { 8'h15, 4'h5 }: pattern = 8'b01101100; 
    { 8'h15, 4'h6 }: pattern = 8'b11000110; 
    { 8'h15, 4'h7 }: pattern = 8'b11000110; 
    { 8'h15, 4'h8 }: pattern = 8'b01101100; 
    { 8'h15, 4'h9 }: pattern = 8'b00111000; 
    { 8'h15, 4'ha }: pattern = 8'b00001100; 
    { 8'h15, 4'hb }: pattern = 8'b11000110; 
    { 8'h15, 4'hc }: pattern = 8'b01111100; 
    { 8'h15, 4'hd }: pattern = 8'b00000000; 
    { 8'h15, 4'he }: pattern = 8'b00000000; 
    { 8'h15, 4'hf }: pattern = 8'b00000000; 

    { 8'h16, 4'h0 }: pattern = 8'b00000000; 
    { 8'h16, 4'h1 }: pattern = 8'b00000000; 
    { 8'h16, 4'h2 }: pattern = 8'b00000000; 
    { 8'h16, 4'h3 }: pattern = 8'b00000000; 
    { 8'h16, 4'h4 }: pattern = 8'b00000000; 
    { 8'h16, 4'h5 }: pattern = 8'b00000000; 
    { 8'h16, 4'h6 }: pattern = 8'b00000000; 
    { 8'h16, 4'h7 }: pattern = 8'b00000000; 
    { 8'h16, 4'h8 }: pattern = 8'b11111110; 
    { 8'h16, 4'h9 }: pattern = 8'b11111110; 
    { 8'h16, 4'ha }: pattern = 8'b11111110; 
    { 8'h16, 4'hb }: pattern = 8'b11111110; 
    { 8'h16, 4'hc }: pattern = 8'b00000000; 
    { 8'h16, 4'hd }: pattern = 8'b00000000; 
    { 8'h16, 4'he }: pattern = 8'b00000000; 
    { 8'h16, 4'hf }: pattern = 8'b00000000; 

    { 8'h17, 4'h0 }: pattern = 8'b00000000; 
    { 8'h17, 4'h1 }: pattern = 8'b00000000; 
    { 8'h17, 4'h2 }: pattern = 8'b00011000; 
    { 8'h17, 4'h3 }: pattern = 8'b00111100; 
    { 8'h17, 4'h4 }: pattern = 8'b01111110; 
    { 8'h17, 4'h5 }: pattern = 8'b00011000; 
    { 8'h17, 4'h6 }: pattern = 8'b00011000; 
    { 8'h17, 4'h7 }: pattern = 8'b00011000; 
    { 8'h17, 4'h8 }: pattern = 8'b01111110; 
    { 8'h17, 4'h9 }: pattern = 8'b00111100; 
    { 8'h17, 4'ha }: pattern = 8'b00011000; 
    { 8'h17, 4'hb }: pattern = 8'b01111110; 
    { 8'h17, 4'hc }: pattern = 8'b00000000; 
    { 8'h17, 4'hd }: pattern = 8'b00000000; 
    { 8'h17, 4'he }: pattern = 8'b00000000; 
    { 8'h17, 4'hf }: pattern = 8'b00000000; 

    { 8'h18, 4'h0 }: pattern = 8'b00000000; 
    { 8'h18, 4'h1 }: pattern = 8'b00000000; 
    { 8'h18, 4'h2 }: pattern = 8'b00011000; 
    { 8'h18, 4'h3 }: pattern = 8'b00111100; 
    { 8'h18, 4'h4 }: pattern = 8'b01111110; 
    { 8'h18, 4'h5 }: pattern = 8'b00011000; 
    { 8'h18, 4'h6 }: pattern = 8'b00011000; 
    { 8'h18, 4'h7 }: pattern = 8'b00011000; 
    { 8'h18, 4'h8 }: pattern = 8'b00011000; 
    { 8'h18, 4'h9 }: pattern = 8'b00011000; 
    { 8'h18, 4'ha }: pattern = 8'b00011000; 
    { 8'h18, 4'hb }: pattern = 8'b00011000; 
    { 8'h18, 4'hc }: pattern = 8'b00000000; 
    { 8'h18, 4'hd }: pattern = 8'b00000000; 
    { 8'h18, 4'he }: pattern = 8'b00000000; 
    { 8'h18, 4'hf }: pattern = 8'b00000000; 

    { 8'h19, 4'h0 }: pattern = 8'b00000000; 
    { 8'h19, 4'h1 }: pattern = 8'b00000000; 
    { 8'h19, 4'h2 }: pattern = 8'b00011000; 
    { 8'h19, 4'h3 }: pattern = 8'b00011000; 
    { 8'h19, 4'h4 }: pattern = 8'b00011000; 
    { 8'h19, 4'h5 }: pattern = 8'b00011000; 
    { 8'h19, 4'h6 }: pattern = 8'b00011000; 
    { 8'h19, 4'h7 }: pattern = 8'b00011000; 
    { 8'h19, 4'h8 }: pattern = 8'b00011000; 
    { 8'h19, 4'h9 }: pattern = 8'b01111110; 
    { 8'h19, 4'ha }: pattern = 8'b00111100; 
    { 8'h19, 4'hb }: pattern = 8'b00011000; 
    { 8'h19, 4'hc }: pattern = 8'b00000000; 
    { 8'h19, 4'hd }: pattern = 8'b00000000; 
    { 8'h19, 4'he }: pattern = 8'b00000000; 
    { 8'h19, 4'hf }: pattern = 8'b00000000; 

    { 8'h1a, 4'h0 }: pattern = 8'b00000000; 
    { 8'h1a, 4'h1 }: pattern = 8'b00000000; 
    { 8'h1a, 4'h2 }: pattern = 8'b00000000; 
    { 8'h1a, 4'h3 }: pattern = 8'b00000000; 
    { 8'h1a, 4'h4 }: pattern = 8'b00000000; 
    { 8'h1a, 4'h5 }: pattern = 8'b00011000; 
    { 8'h1a, 4'h6 }: pattern = 8'b00001100; 
    { 8'h1a, 4'h7 }: pattern = 8'b11111110; 
    { 8'h1a, 4'h8 }: pattern = 8'b00001100; 
    { 8'h1a, 4'h9 }: pattern = 8'b00011000; 
    { 8'h1a, 4'ha }: pattern = 8'b00000000; 
    { 8'h1a, 4'hb }: pattern = 8'b00000000; 
    { 8'h1a, 4'hc }: pattern = 8'b00000000; 
    { 8'h1a, 4'hd }: pattern = 8'b00000000; 
    { 8'h1a, 4'he }: pattern = 8'b00000000; 
    { 8'h1a, 4'hf }: pattern = 8'b00000000; 

    { 8'h1b, 4'h0 }: pattern = 8'b00000000; 
    { 8'h1b, 4'h1 }: pattern = 8'b00000000; 
    { 8'h1b, 4'h2 }: pattern = 8'b00000000; 
    { 8'h1b, 4'h3 }: pattern = 8'b00000000; 
    { 8'h1b, 4'h4 }: pattern = 8'b00000000; 
    { 8'h1b, 4'h5 }: pattern = 8'b00110000; 
    { 8'h1b, 4'h6 }: pattern = 8'b01100000; 
    { 8'h1b, 4'h7 }: pattern = 8'b11111110; 
    { 8'h1b, 4'h8 }: pattern = 8'b01100000; 
    { 8'h1b, 4'h9 }: pattern = 8'b00110000; 
    { 8'h1b, 4'ha }: pattern = 8'b00000000; 
    { 8'h1b, 4'hb }: pattern = 8'b00000000; 
    { 8'h1b, 4'hc }: pattern = 8'b00000000; 
    { 8'h1b, 4'hd }: pattern = 8'b00000000; 
    { 8'h1b, 4'he }: pattern = 8'b00000000; 
    { 8'h1b, 4'hf }: pattern = 8'b00000000; 

    { 8'h1c, 4'h0 }: pattern = 8'b00000000; 
    { 8'h1c, 4'h1 }: pattern = 8'b00000000; 
    { 8'h1c, 4'h2 }: pattern = 8'b00000000; 
    { 8'h1c, 4'h3 }: pattern = 8'b00000000; 
    { 8'h1c, 4'h4 }: pattern = 8'b00000000; 
    { 8'h1c, 4'h5 }: pattern = 8'b00000000; 
    { 8'h1c, 4'h6 }: pattern = 8'b11000000; 
    { 8'h1c, 4'h7 }: pattern = 8'b11000000; 
    { 8'h1c, 4'h8 }: pattern = 8'b11000000; 
    { 8'h1c, 4'h9 }: pattern = 8'b11111110; 
    { 8'h1c, 4'ha }: pattern = 8'b00000000; 
    { 8'h1c, 4'hb }: pattern = 8'b00000000; 
    { 8'h1c, 4'hc }: pattern = 8'b00000000; 
    { 8'h1c, 4'hd }: pattern = 8'b00000000; 
    { 8'h1c, 4'he }: pattern = 8'b00000000; 
    { 8'h1c, 4'hf }: pattern = 8'b00000000; 

    { 8'h1d, 4'h0 }: pattern = 8'b00000000; 
    { 8'h1d, 4'h1 }: pattern = 8'b00000000; 
    { 8'h1d, 4'h2 }: pattern = 8'b00000000; 
    { 8'h1d, 4'h3 }: pattern = 8'b00000000; 
    { 8'h1d, 4'h4 }: pattern = 8'b00000000; 
    { 8'h1d, 4'h5 }: pattern = 8'b00101000; 
    { 8'h1d, 4'h6 }: pattern = 8'b01101100; 
    { 8'h1d, 4'h7 }: pattern = 8'b11111110; 
    { 8'h1d, 4'h8 }: pattern = 8'b01101100; 
    { 8'h1d, 4'h9 }: pattern = 8'b00101000; 
    { 8'h1d, 4'ha }: pattern = 8'b00000000; 
    { 8'h1d, 4'hb }: pattern = 8'b00000000; 
    { 8'h1d, 4'hc }: pattern = 8'b00000000; 
    { 8'h1d, 4'hd }: pattern = 8'b00000000; 
    { 8'h1d, 4'he }: pattern = 8'b00000000; 
    { 8'h1d, 4'hf }: pattern = 8'b00000000; 

    { 8'h1e, 4'h0 }: pattern = 8'b00000000; 
    { 8'h1e, 4'h1 }: pattern = 8'b00000000; 
    { 8'h1e, 4'h2 }: pattern = 8'b00000000; 
    { 8'h1e, 4'h3 }: pattern = 8'b00000000; 
    { 8'h1e, 4'h4 }: pattern = 8'b00010000; 
    { 8'h1e, 4'h5 }: pattern = 8'b00111000; 
    { 8'h1e, 4'h6 }: pattern = 8'b00111000; 
    { 8'h1e, 4'h7 }: pattern = 8'b01111100; 
    { 8'h1e, 4'h8 }: pattern = 8'b01111100; 
    { 8'h1e, 4'h9 }: pattern = 8'b11111110; 
    { 8'h1e, 4'ha }: pattern = 8'b11111110; 
    { 8'h1e, 4'hb }: pattern = 8'b00000000; 
    { 8'h1e, 4'hc }: pattern = 8'b00000000; 
    { 8'h1e, 4'hd }: pattern = 8'b00000000; 
    { 8'h1e, 4'he }: pattern = 8'b00000000; 
    { 8'h1e, 4'hf }: pattern = 8'b00000000; 

    { 8'h1f, 4'h0 }: pattern = 8'b00000000; 
    { 8'h1f, 4'h1 }: pattern = 8'b00000000; 
    { 8'h1f, 4'h2 }: pattern = 8'b00000000; 
    { 8'h1f, 4'h3 }: pattern = 8'b00000000; 
    { 8'h1f, 4'h4 }: pattern = 8'b11111110; 
    { 8'h1f, 4'h5 }: pattern = 8'b11111110; 
    { 8'h1f, 4'h6 }: pattern = 8'b01111100; 
    { 8'h1f, 4'h7 }: pattern = 8'b01111100; 
    { 8'h1f, 4'h8 }: pattern = 8'b00111000; 
    { 8'h1f, 4'h9 }: pattern = 8'b00111000; 
    { 8'h1f, 4'ha }: pattern = 8'b00010000; 
    { 8'h1f, 4'hb }: pattern = 8'b00000000; 
    { 8'h1f, 4'hc }: pattern = 8'b00000000; 
    { 8'h1f, 4'hd }: pattern = 8'b00000000; 
    { 8'h1f, 4'he }: pattern = 8'b00000000; 
    { 8'h1f, 4'hf }: pattern = 8'b00000000; 

    { 8'h20, 4'h0 }: pattern = 8'b00000000; 
    { 8'h20, 4'h1 }: pattern = 8'b00000000; 
    { 8'h20, 4'h2 }: pattern = 8'b00000000; 
    { 8'h20, 4'h3 }: pattern = 8'b00000000; 
    { 8'h20, 4'h4 }: pattern = 8'b00000000; 
    { 8'h20, 4'h5 }: pattern = 8'b00000000; 
    { 8'h20, 4'h6 }: pattern = 8'b00000000; 
    { 8'h20, 4'h7 }: pattern = 8'b00000000; 
    { 8'h20, 4'h8 }: pattern = 8'b00000000; 
    { 8'h20, 4'h9 }: pattern = 8'b00000000; 
    { 8'h20, 4'ha }: pattern = 8'b00000000; 
    { 8'h20, 4'hb }: pattern = 8'b00000000; 
    { 8'h20, 4'hc }: pattern = 8'b00000000; 
    { 8'h20, 4'hd }: pattern = 8'b00000000; 
    { 8'h20, 4'he }: pattern = 8'b00000000; 
    { 8'h20, 4'hf }: pattern = 8'b00000000; 

    { 8'h21, 4'h0 }: pattern = 8'b00000000; 
    { 8'h21, 4'h1 }: pattern = 8'b00000000; 
    { 8'h21, 4'h2 }: pattern = 8'b00011000; 
    { 8'h21, 4'h3 }: pattern = 8'b00111100; 
    { 8'h21, 4'h4 }: pattern = 8'b00111100; 
    { 8'h21, 4'h5 }: pattern = 8'b00111100; 
    { 8'h21, 4'h6 }: pattern = 8'b00011000; 
    { 8'h21, 4'h7 }: pattern = 8'b00011000; 
    { 8'h21, 4'h8 }: pattern = 8'b00011000; 
    { 8'h21, 4'h9 }: pattern = 8'b00000000; 
    { 8'h21, 4'ha }: pattern = 8'b00011000; 
    { 8'h21, 4'hb }: pattern = 8'b00011000; 
    { 8'h21, 4'hc }: pattern = 8'b00000000; 
    { 8'h21, 4'hd }: pattern = 8'b00000000; 
    { 8'h21, 4'he }: pattern = 8'b00000000; 
    { 8'h21, 4'hf }: pattern = 8'b00000000; 

    { 8'h22, 4'h0 }: pattern = 8'b00000000; 
    { 8'h22, 4'h1 }: pattern = 8'b01100110; 
    { 8'h22, 4'h2 }: pattern = 8'b01100110; 
    { 8'h22, 4'h3 }: pattern = 8'b01100110; 
    { 8'h22, 4'h4 }: pattern = 8'b00100100; 
    { 8'h22, 4'h5 }: pattern = 8'b00000000; 
    { 8'h22, 4'h6 }: pattern = 8'b00000000; 
    { 8'h22, 4'h7 }: pattern = 8'b00000000; 
    { 8'h22, 4'h8 }: pattern = 8'b00000000; 
    { 8'h22, 4'h9 }: pattern = 8'b00000000; 
    { 8'h22, 4'ha }: pattern = 8'b00000000; 
    { 8'h22, 4'hb }: pattern = 8'b00000000; 
    { 8'h22, 4'hc }: pattern = 8'b00000000; 
    { 8'h22, 4'hd }: pattern = 8'b00000000; 
    { 8'h22, 4'he }: pattern = 8'b00000000; 
    { 8'h22, 4'hf }: pattern = 8'b00000000; 

    { 8'h23, 4'h0 }: pattern = 8'b00000000; 
    { 8'h23, 4'h1 }: pattern = 8'b00000000; 
    { 8'h23, 4'h2 }: pattern = 8'b00000000; 
    { 8'h23, 4'h3 }: pattern = 8'b01101100; 
    { 8'h23, 4'h4 }: pattern = 8'b01101100; 
    { 8'h23, 4'h5 }: pattern = 8'b11111110; 
    { 8'h23, 4'h6 }: pattern = 8'b01101100; 
    { 8'h23, 4'h7 }: pattern = 8'b01101100; 
    { 8'h23, 4'h8 }: pattern = 8'b01101100; 
    { 8'h23, 4'h9 }: pattern = 8'b11111110; 
    { 8'h23, 4'ha }: pattern = 8'b01101100; 
    { 8'h23, 4'hb }: pattern = 8'b01101100; 
    { 8'h23, 4'hc }: pattern = 8'b00000000; 
    { 8'h23, 4'hd }: pattern = 8'b00000000; 
    { 8'h23, 4'he }: pattern = 8'b00000000; 
    { 8'h23, 4'hf }: pattern = 8'b00000000; 

    { 8'h24, 4'h0 }: pattern = 8'b00011000; 
    { 8'h24, 4'h1 }: pattern = 8'b00011000; 
    { 8'h24, 4'h2 }: pattern = 8'b01111100; 
    { 8'h24, 4'h3 }: pattern = 8'b11000110; 
    { 8'h24, 4'h4 }: pattern = 8'b11000010; 
    { 8'h24, 4'h5 }: pattern = 8'b11000000; 
    { 8'h24, 4'h6 }: pattern = 8'b01111100; 
    { 8'h24, 4'h7 }: pattern = 8'b00000110; 
    { 8'h24, 4'h8 }: pattern = 8'b00000110; 
    { 8'h24, 4'h9 }: pattern = 8'b10000110; 
    { 8'h24, 4'ha }: pattern = 8'b11000110; 
    { 8'h24, 4'hb }: pattern = 8'b01111100; 
    { 8'h24, 4'hc }: pattern = 8'b00011000; 
    { 8'h24, 4'hd }: pattern = 8'b00011000; 
    { 8'h24, 4'he }: pattern = 8'b00000000; 
    { 8'h24, 4'hf }: pattern = 8'b00000000; 

    { 8'h25, 4'h0 }: pattern = 8'b00000000; 
    { 8'h25, 4'h1 }: pattern = 8'b00000000; 
    { 8'h25, 4'h2 }: pattern = 8'b00000000; 
    { 8'h25, 4'h3 }: pattern = 8'b00000000; 
    { 8'h25, 4'h4 }: pattern = 8'b11000010; 
    { 8'h25, 4'h5 }: pattern = 8'b11000110; 
    { 8'h25, 4'h6 }: pattern = 8'b00001100; 
    { 8'h25, 4'h7 }: pattern = 8'b00011000; 
    { 8'h25, 4'h8 }: pattern = 8'b00110000; 
    { 8'h25, 4'h9 }: pattern = 8'b01100000; 
    { 8'h25, 4'ha }: pattern = 8'b11000110; 
    { 8'h25, 4'hb }: pattern = 8'b10000110; 
    { 8'h25, 4'hc }: pattern = 8'b00000000; 
    { 8'h25, 4'hd }: pattern = 8'b00000000; 
    { 8'h25, 4'he }: pattern = 8'b00000000; 
    { 8'h25, 4'hf }: pattern = 8'b00000000; 

    { 8'h26, 4'h0 }: pattern = 8'b00000000; 
    { 8'h26, 4'h1 }: pattern = 8'b00000000; 
    { 8'h26, 4'h2 }: pattern = 8'b00111000; 
    { 8'h26, 4'h3 }: pattern = 8'b01101100; 
    { 8'h26, 4'h4 }: pattern = 8'b01101100; 
    { 8'h26, 4'h5 }: pattern = 8'b00111000; 
    { 8'h26, 4'h6 }: pattern = 8'b01110110; 
    { 8'h26, 4'h7 }: pattern = 8'b11011100; 
    { 8'h26, 4'h8 }: pattern = 8'b11001100; 
    { 8'h26, 4'h9 }: pattern = 8'b11001100; 
    { 8'h26, 4'ha }: pattern = 8'b11001100; 
    { 8'h26, 4'hb }: pattern = 8'b01110110; 
    { 8'h26, 4'hc }: pattern = 8'b00000000; 
    { 8'h26, 4'hd }: pattern = 8'b00000000; 
    { 8'h26, 4'he }: pattern = 8'b00000000; 
    { 8'h26, 4'hf }: pattern = 8'b00000000; 

    { 8'h27, 4'h0 }: pattern = 8'b00000000; 
    { 8'h27, 4'h1 }: pattern = 8'b00110000; 
    { 8'h27, 4'h2 }: pattern = 8'b00110000; 
    { 8'h27, 4'h3 }: pattern = 8'b00110000; 
    { 8'h27, 4'h4 }: pattern = 8'b01100000; 
    { 8'h27, 4'h5 }: pattern = 8'b00000000; 
    { 8'h27, 4'h6 }: pattern = 8'b00000000; 
    { 8'h27, 4'h7 }: pattern = 8'b00000000; 
    { 8'h27, 4'h8 }: pattern = 8'b00000000; 
    { 8'h27, 4'h9 }: pattern = 8'b00000000; 
    { 8'h27, 4'ha }: pattern = 8'b00000000; 
    { 8'h27, 4'hb }: pattern = 8'b00000000; 
    { 8'h27, 4'hc }: pattern = 8'b00000000; 
    { 8'h27, 4'hd }: pattern = 8'b00000000; 
    { 8'h27, 4'he }: pattern = 8'b00000000; 
    { 8'h27, 4'hf }: pattern = 8'b00000000; 

    { 8'h28, 4'h0 }: pattern = 8'b00000000; 
    { 8'h28, 4'h1 }: pattern = 8'b00000000; 
    { 8'h28, 4'h2 }: pattern = 8'b00001100; 
    { 8'h28, 4'h3 }: pattern = 8'b00011000; 
    { 8'h28, 4'h4 }: pattern = 8'b00110000; 
    { 8'h28, 4'h5 }: pattern = 8'b00110000; 
    { 8'h28, 4'h6 }: pattern = 8'b00110000; 
    { 8'h28, 4'h7 }: pattern = 8'b00110000; 
    { 8'h28, 4'h8 }: pattern = 8'b00110000; 
    { 8'h28, 4'h9 }: pattern = 8'b00110000; 
    { 8'h28, 4'ha }: pattern = 8'b00011000; 
    { 8'h28, 4'hb }: pattern = 8'b00001100; 
    { 8'h28, 4'hc }: pattern = 8'b00000000; 
    { 8'h28, 4'hd }: pattern = 8'b00000000; 
    { 8'h28, 4'he }: pattern = 8'b00000000; 
    { 8'h28, 4'hf }: pattern = 8'b00000000; 

    { 8'h29, 4'h0 }: pattern = 8'b00000000; 
    { 8'h29, 4'h1 }: pattern = 8'b00000000; 
    { 8'h29, 4'h2 }: pattern = 8'b00110000; 
    { 8'h29, 4'h3 }: pattern = 8'b00011000; 
    { 8'h29, 4'h4 }: pattern = 8'b00001100; 
    { 8'h29, 4'h5 }: pattern = 8'b00001100; 
    { 8'h29, 4'h6 }: pattern = 8'b00001100; 
    { 8'h29, 4'h7 }: pattern = 8'b00001100; 
    { 8'h29, 4'h8 }: pattern = 8'b00001100; 
    { 8'h29, 4'h9 }: pattern = 8'b00001100; 
    { 8'h29, 4'ha }: pattern = 8'b00011000; 
    { 8'h29, 4'hb }: pattern = 8'b00110000; 
    { 8'h29, 4'hc }: pattern = 8'b00000000; 
    { 8'h29, 4'hd }: pattern = 8'b00000000; 
    { 8'h29, 4'he }: pattern = 8'b00000000; 
    { 8'h29, 4'hf }: pattern = 8'b00000000; 

    { 8'h2a, 4'h0 }: pattern = 8'b00000000; 
    { 8'h2a, 4'h1 }: pattern = 8'b00000000; 
    { 8'h2a, 4'h2 }: pattern = 8'b00000000; 
    { 8'h2a, 4'h3 }: pattern = 8'b00000000; 
    { 8'h2a, 4'h4 }: pattern = 8'b00000000; 
    { 8'h2a, 4'h5 }: pattern = 8'b01100110; 
    { 8'h2a, 4'h6 }: pattern = 8'b00111100; 
    { 8'h2a, 4'h7 }: pattern = 8'b11111111; 
    { 8'h2a, 4'h8 }: pattern = 8'b00111100; 
    { 8'h2a, 4'h9 }: pattern = 8'b01100110; 
    { 8'h2a, 4'ha }: pattern = 8'b00000000; 
    { 8'h2a, 4'hb }: pattern = 8'b00000000; 
    { 8'h2a, 4'hc }: pattern = 8'b00000000; 
    { 8'h2a, 4'hd }: pattern = 8'b00000000; 
    { 8'h2a, 4'he }: pattern = 8'b00000000; 
    { 8'h2a, 4'hf }: pattern = 8'b00000000; 

    { 8'h2b, 4'h0 }: pattern = 8'b00000000; 
    { 8'h2b, 4'h1 }: pattern = 8'b00000000; 
    { 8'h2b, 4'h2 }: pattern = 8'b00000000; 
    { 8'h2b, 4'h3 }: pattern = 8'b00000000; 
    { 8'h2b, 4'h4 }: pattern = 8'b00000000; 
    { 8'h2b, 4'h5 }: pattern = 8'b00011000; 
    { 8'h2b, 4'h6 }: pattern = 8'b00011000; 
    { 8'h2b, 4'h7 }: pattern = 8'b01111110; 
    { 8'h2b, 4'h8 }: pattern = 8'b00011000; 
    { 8'h2b, 4'h9 }: pattern = 8'b00011000; 
    { 8'h2b, 4'ha }: pattern = 8'b00000000; 
    { 8'h2b, 4'hb }: pattern = 8'b00000000; 
    { 8'h2b, 4'hc }: pattern = 8'b00000000; 
    { 8'h2b, 4'hd }: pattern = 8'b00000000; 
    { 8'h2b, 4'he }: pattern = 8'b00000000; 
    { 8'h2b, 4'hf }: pattern = 8'b00000000; 

    { 8'h2c, 4'h0 }: pattern = 8'b00000000; 
    { 8'h2c, 4'h1 }: pattern = 8'b00000000; 
    { 8'h2c, 4'h2 }: pattern = 8'b00000000; 
    { 8'h2c, 4'h3 }: pattern = 8'b00000000; 
    { 8'h2c, 4'h4 }: pattern = 8'b00000000; 
    { 8'h2c, 4'h5 }: pattern = 8'b00000000; 
    { 8'h2c, 4'h6 }: pattern = 8'b00000000; 
    { 8'h2c, 4'h7 }: pattern = 8'b00000000; 
    { 8'h2c, 4'h8 }: pattern = 8'b00000000; 
    { 8'h2c, 4'h9 }: pattern = 8'b00011000; 
    { 8'h2c, 4'ha }: pattern = 8'b00011000; 
    { 8'h2c, 4'hb }: pattern = 8'b00011000; 
    { 8'h2c, 4'hc }: pattern = 8'b00110000; 
    { 8'h2c, 4'hd }: pattern = 8'b00000000; 
    { 8'h2c, 4'he }: pattern = 8'b00000000; 
    { 8'h2c, 4'hf }: pattern = 8'b00000000; 

    { 8'h2d, 4'h0 }: pattern = 8'b00000000; 
    { 8'h2d, 4'h1 }: pattern = 8'b00000000; 
    { 8'h2d, 4'h2 }: pattern = 8'b00000000; 
    { 8'h2d, 4'h3 }: pattern = 8'b00000000; 
    { 8'h2d, 4'h4 }: pattern = 8'b00000000; 
    { 8'h2d, 4'h5 }: pattern = 8'b00000000; 
    { 8'h2d, 4'h6 }: pattern = 8'b00000000; 
    { 8'h2d, 4'h7 }: pattern = 8'b11111110; 
    { 8'h2d, 4'h8 }: pattern = 8'b00000000; 
    { 8'h2d, 4'h9 }: pattern = 8'b00000000; 
    { 8'h2d, 4'ha }: pattern = 8'b00000000; 
    { 8'h2d, 4'hb }: pattern = 8'b00000000; 
    { 8'h2d, 4'hc }: pattern = 8'b00000000; 
    { 8'h2d, 4'hd }: pattern = 8'b00000000; 
    { 8'h2d, 4'he }: pattern = 8'b00000000; 
    { 8'h2d, 4'hf }: pattern = 8'b00000000; 

    { 8'h2e, 4'h0 }: pattern = 8'b00000000; 
    { 8'h2e, 4'h1 }: pattern = 8'b00000000; 
    { 8'h2e, 4'h2 }: pattern = 8'b00000000; 
    { 8'h2e, 4'h3 }: pattern = 8'b00000000; 
    { 8'h2e, 4'h4 }: pattern = 8'b00000000; 
    { 8'h2e, 4'h5 }: pattern = 8'b00000000; 
    { 8'h2e, 4'h6 }: pattern = 8'b00000000; 
    { 8'h2e, 4'h7 }: pattern = 8'b00000000; 
    { 8'h2e, 4'h8 }: pattern = 8'b00000000; 
    { 8'h2e, 4'h9 }: pattern = 8'b00000000; 
    { 8'h2e, 4'ha }: pattern = 8'b00011000; 
    { 8'h2e, 4'hb }: pattern = 8'b00011000; 
    { 8'h2e, 4'hc }: pattern = 8'b00000000; 
    { 8'h2e, 4'hd }: pattern = 8'b00000000; 
    { 8'h2e, 4'he }: pattern = 8'b00000000; 
    { 8'h2e, 4'hf }: pattern = 8'b00000000; 

    { 8'h2f, 4'h0 }: pattern = 8'b00000000; 
    { 8'h2f, 4'h1 }: pattern = 8'b00000000; 
    { 8'h2f, 4'h2 }: pattern = 8'b00000000; 
    { 8'h2f, 4'h3 }: pattern = 8'b00000000; 
    { 8'h2f, 4'h4 }: pattern = 8'b00000010; 
    { 8'h2f, 4'h5 }: pattern = 8'b00000110; 
    { 8'h2f, 4'h6 }: pattern = 8'b00001100; 
    { 8'h2f, 4'h7 }: pattern = 8'b00011000; 
    { 8'h2f, 4'h8 }: pattern = 8'b00110000; 
    { 8'h2f, 4'h9 }: pattern = 8'b01100000; 
    { 8'h2f, 4'ha }: pattern = 8'b11000000; 
    { 8'h2f, 4'hb }: pattern = 8'b10000000; 
    { 8'h2f, 4'hc }: pattern = 8'b00000000; 
    { 8'h2f, 4'hd }: pattern = 8'b00000000; 
    { 8'h2f, 4'he }: pattern = 8'b00000000; 
    { 8'h2f, 4'hf }: pattern = 8'b00000000; 

    { 8'h30, 4'h0 }: pattern = 8'b00000000; 
    { 8'h30, 4'h1 }: pattern = 8'b00000000; 
    { 8'h30, 4'h2 }: pattern = 8'b00111000; 
    { 8'h30, 4'h3 }: pattern = 8'b01101100; 
    { 8'h30, 4'h4 }: pattern = 8'b11000110; 
    { 8'h30, 4'h5 }: pattern = 8'b11000110; 
    { 8'h30, 4'h6 }: pattern = 8'b11010110; 
    { 8'h30, 4'h7 }: pattern = 8'b11010110; 
    { 8'h30, 4'h8 }: pattern = 8'b11000110; 
    { 8'h30, 4'h9 }: pattern = 8'b11000110; 
    { 8'h30, 4'ha }: pattern = 8'b01101100; 
    { 8'h30, 4'hb }: pattern = 8'b00111000; 
    { 8'h30, 4'hc }: pattern = 8'b00000000; 
    { 8'h30, 4'hd }: pattern = 8'b00000000; 
    { 8'h30, 4'he }: pattern = 8'b00000000; 
    { 8'h30, 4'hf }: pattern = 8'b00000000; 

    { 8'h31, 4'h0 }: pattern = 8'b00000000; 
    { 8'h31, 4'h1 }: pattern = 8'b00000000; 
    { 8'h31, 4'h2 }: pattern = 8'b00011000; 
    { 8'h31, 4'h3 }: pattern = 8'b00111000; 
    { 8'h31, 4'h4 }: pattern = 8'b01111000; 
    { 8'h31, 4'h5 }: pattern = 8'b00011000; 
    { 8'h31, 4'h6 }: pattern = 8'b00011000; 
    { 8'h31, 4'h7 }: pattern = 8'b00011000; 
    { 8'h31, 4'h8 }: pattern = 8'b00011000; 
    { 8'h31, 4'h9 }: pattern = 8'b00011000; 
    { 8'h31, 4'ha }: pattern = 8'b00011000; 
    { 8'h31, 4'hb }: pattern = 8'b01111110; 
    { 8'h31, 4'hc }: pattern = 8'b00000000; 
    { 8'h31, 4'hd }: pattern = 8'b00000000; 
    { 8'h31, 4'he }: pattern = 8'b00000000; 
    { 8'h31, 4'hf }: pattern = 8'b00000000; 

    { 8'h32, 4'h0 }: pattern = 8'b00000000; 
    { 8'h32, 4'h1 }: pattern = 8'b00000000; 
    { 8'h32, 4'h2 }: pattern = 8'b01111100; 
    { 8'h32, 4'h3 }: pattern = 8'b11000110; 
    { 8'h32, 4'h4 }: pattern = 8'b00000110; 
    { 8'h32, 4'h5 }: pattern = 8'b00001100; 
    { 8'h32, 4'h6 }: pattern = 8'b00011000; 
    { 8'h32, 4'h7 }: pattern = 8'b00110000; 
    { 8'h32, 4'h8 }: pattern = 8'b01100000; 
    { 8'h32, 4'h9 }: pattern = 8'b11000000; 
    { 8'h32, 4'ha }: pattern = 8'b11000110; 
    { 8'h32, 4'hb }: pattern = 8'b11111110; 
    { 8'h32, 4'hc }: pattern = 8'b00000000; 
    { 8'h32, 4'hd }: pattern = 8'b00000000; 
    { 8'h32, 4'he }: pattern = 8'b00000000; 
    { 8'h32, 4'hf }: pattern = 8'b00000000; 

    { 8'h33, 4'h0 }: pattern = 8'b00000000; 
    { 8'h33, 4'h1 }: pattern = 8'b00000000; 
    { 8'h33, 4'h2 }: pattern = 8'b01111100; 
    { 8'h33, 4'h3 }: pattern = 8'b11000110; 
    { 8'h33, 4'h4 }: pattern = 8'b00000110; 
    { 8'h33, 4'h5 }: pattern = 8'b00000110; 
    { 8'h33, 4'h6 }: pattern = 8'b00111100; 
    { 8'h33, 4'h7 }: pattern = 8'b00000110; 
    { 8'h33, 4'h8 }: pattern = 8'b00000110; 
    { 8'h33, 4'h9 }: pattern = 8'b00000110; 
    { 8'h33, 4'ha }: pattern = 8'b11000110; 
    { 8'h33, 4'hb }: pattern = 8'b01111100; 
    { 8'h33, 4'hc }: pattern = 8'b00000000; 
    { 8'h33, 4'hd }: pattern = 8'b00000000; 
    { 8'h33, 4'he }: pattern = 8'b00000000; 
    { 8'h33, 4'hf }: pattern = 8'b00000000; 

    { 8'h34, 4'h0 }: pattern = 8'b00000000; 
    { 8'h34, 4'h1 }: pattern = 8'b00000000; 
    { 8'h34, 4'h2 }: pattern = 8'b00001100; 
    { 8'h34, 4'h3 }: pattern = 8'b00011100; 
    { 8'h34, 4'h4 }: pattern = 8'b00111100; 
    { 8'h34, 4'h5 }: pattern = 8'b01101100; 
    { 8'h34, 4'h6 }: pattern = 8'b11001100; 
    { 8'h34, 4'h7 }: pattern = 8'b11111110; 
    { 8'h34, 4'h8 }: pattern = 8'b00001100; 
    { 8'h34, 4'h9 }: pattern = 8'b00001100; 
    { 8'h34, 4'ha }: pattern = 8'b00001100; 
    { 8'h34, 4'hb }: pattern = 8'b00011110; 
    { 8'h34, 4'hc }: pattern = 8'b00000000; 
    { 8'h34, 4'hd }: pattern = 8'b00000000; 
    { 8'h34, 4'he }: pattern = 8'b00000000; 
    { 8'h34, 4'hf }: pattern = 8'b00000000; 

    { 8'h35, 4'h0 }: pattern = 8'b00000000; 
    { 8'h35, 4'h1 }: pattern = 8'b00000000; 
    { 8'h35, 4'h2 }: pattern = 8'b11111110; 
    { 8'h35, 4'h3 }: pattern = 8'b11000000; 
    { 8'h35, 4'h4 }: pattern = 8'b11000000; 
    { 8'h35, 4'h5 }: pattern = 8'b11000000; 
    { 8'h35, 4'h6 }: pattern = 8'b11111100; 
    { 8'h35, 4'h7 }: pattern = 8'b00000110; 
    { 8'h35, 4'h8 }: pattern = 8'b00000110; 
    { 8'h35, 4'h9 }: pattern = 8'b00000110; 
    { 8'h35, 4'ha }: pattern = 8'b11000110; 
    { 8'h35, 4'hb }: pattern = 8'b01111100; 
    { 8'h35, 4'hc }: pattern = 8'b00000000; 
    { 8'h35, 4'hd }: pattern = 8'b00000000; 
    { 8'h35, 4'he }: pattern = 8'b00000000; 
    { 8'h35, 4'hf }: pattern = 8'b00000000; 

    { 8'h36, 4'h0 }: pattern = 8'b00000000; 
    { 8'h36, 4'h1 }: pattern = 8'b00000000; 
    { 8'h36, 4'h2 }: pattern = 8'b00111000; 
    { 8'h36, 4'h3 }: pattern = 8'b01100000; 
    { 8'h36, 4'h4 }: pattern = 8'b11000000; 
    { 8'h36, 4'h5 }: pattern = 8'b11000000; 
    { 8'h36, 4'h6 }: pattern = 8'b11111100; 
    { 8'h36, 4'h7 }: pattern = 8'b11000110; 
    { 8'h36, 4'h8 }: pattern = 8'b11000110; 
    { 8'h36, 4'h9 }: pattern = 8'b11000110; 
    { 8'h36, 4'ha }: pattern = 8'b11000110; 
    { 8'h36, 4'hb }: pattern = 8'b01111100; 
    { 8'h36, 4'hc }: pattern = 8'b00000000; 
    { 8'h36, 4'hd }: pattern = 8'b00000000; 
    { 8'h36, 4'he }: pattern = 8'b00000000; 
    { 8'h36, 4'hf }: pattern = 8'b00000000; 

    { 8'h37, 4'h0 }: pattern = 8'b00000000; 
    { 8'h37, 4'h1 }: pattern = 8'b00000000; 
    { 8'h37, 4'h2 }: pattern = 8'b11111110; 
    { 8'h37, 4'h3 }: pattern = 8'b11000110; 
    { 8'h37, 4'h4 }: pattern = 8'b00000110; 
    { 8'h37, 4'h5 }: pattern = 8'b00000110; 
    { 8'h37, 4'h6 }: pattern = 8'b00001100; 
    { 8'h37, 4'h7 }: pattern = 8'b00011000; 
    { 8'h37, 4'h8 }: pattern = 8'b00110000; 
    { 8'h37, 4'h9 }: pattern = 8'b00110000; 
    { 8'h37, 4'ha }: pattern = 8'b00110000; 
    { 8'h37, 4'hb }: pattern = 8'b00110000; 
    { 8'h37, 4'hc }: pattern = 8'b00000000; 
    { 8'h37, 4'hd }: pattern = 8'b00000000; 
    { 8'h37, 4'he }: pattern = 8'b00000000; 
    { 8'h37, 4'hf }: pattern = 8'b00000000; 

    { 8'h38, 4'h0 }: pattern = 8'b00000000; 
    { 8'h38, 4'h1 }: pattern = 8'b00000000; 
    { 8'h38, 4'h2 }: pattern = 8'b01111100; 
    { 8'h38, 4'h3 }: pattern = 8'b11000110; 
    { 8'h38, 4'h4 }: pattern = 8'b11000110; 
    { 8'h38, 4'h5 }: pattern = 8'b11000110; 
    { 8'h38, 4'h6 }: pattern = 8'b01111100; 
    { 8'h38, 4'h7 }: pattern = 8'b11000110; 
    { 8'h38, 4'h8 }: pattern = 8'b11000110; 
    { 8'h38, 4'h9 }: pattern = 8'b11000110; 
    { 8'h38, 4'ha }: pattern = 8'b11000110; 
    { 8'h38, 4'hb }: pattern = 8'b01111100; 
    { 8'h38, 4'hc }: pattern = 8'b00000000; 
    { 8'h38, 4'hd }: pattern = 8'b00000000; 
    { 8'h38, 4'he }: pattern = 8'b00000000; 
    { 8'h38, 4'hf }: pattern = 8'b00000000; 

    { 8'h39, 4'h0 }: pattern = 8'b00000000; 
    { 8'h39, 4'h1 }: pattern = 8'b00000000; 
    { 8'h39, 4'h2 }: pattern = 8'b01111100; 
    { 8'h39, 4'h3 }: pattern = 8'b11000110; 
    { 8'h39, 4'h4 }: pattern = 8'b11000110; 
    { 8'h39, 4'h5 }: pattern = 8'b11000110; 
    { 8'h39, 4'h6 }: pattern = 8'b01111110; 
    { 8'h39, 4'h7 }: pattern = 8'b00000110; 
    { 8'h39, 4'h8 }: pattern = 8'b00000110; 
    { 8'h39, 4'h9 }: pattern = 8'b00000110; 
    { 8'h39, 4'ha }: pattern = 8'b00001100; 
    { 8'h39, 4'hb }: pattern = 8'b01111000; 
    { 8'h39, 4'hc }: pattern = 8'b00000000; 
    { 8'h39, 4'hd }: pattern = 8'b00000000; 
    { 8'h39, 4'he }: pattern = 8'b00000000; 
    { 8'h39, 4'hf }: pattern = 8'b00000000; 

    { 8'h3a, 4'h0 }: pattern = 8'b00000000; 
    { 8'h3a, 4'h1 }: pattern = 8'b00000000; 
    { 8'h3a, 4'h2 }: pattern = 8'b00000000; 
    { 8'h3a, 4'h3 }: pattern = 8'b00000000; 
    { 8'h3a, 4'h4 }: pattern = 8'b00011000; 
    { 8'h3a, 4'h5 }: pattern = 8'b00011000; 
    { 8'h3a, 4'h6 }: pattern = 8'b00000000; 
    { 8'h3a, 4'h7 }: pattern = 8'b00000000; 
    { 8'h3a, 4'h8 }: pattern = 8'b00000000; 
    { 8'h3a, 4'h9 }: pattern = 8'b00011000; 
    { 8'h3a, 4'ha }: pattern = 8'b00011000; 
    { 8'h3a, 4'hb }: pattern = 8'b00000000; 
    { 8'h3a, 4'hc }: pattern = 8'b00000000; 
    { 8'h3a, 4'hd }: pattern = 8'b00000000; 
    { 8'h3a, 4'he }: pattern = 8'b00000000; 
    { 8'h3a, 4'hf }: pattern = 8'b00000000; 

    { 8'h3b, 4'h0 }: pattern = 8'b00000000; 
    { 8'h3b, 4'h1 }: pattern = 8'b00000000; 
    { 8'h3b, 4'h2 }: pattern = 8'b00000000; 
    { 8'h3b, 4'h3 }: pattern = 8'b00000000; 
    { 8'h3b, 4'h4 }: pattern = 8'b00011000; 
    { 8'h3b, 4'h5 }: pattern = 8'b00011000; 
    { 8'h3b, 4'h6 }: pattern = 8'b00000000; 
    { 8'h3b, 4'h7 }: pattern = 8'b00000000; 
    { 8'h3b, 4'h8 }: pattern = 8'b00000000; 
    { 8'h3b, 4'h9 }: pattern = 8'b00011000; 
    { 8'h3b, 4'ha }: pattern = 8'b00011000; 
    { 8'h3b, 4'hb }: pattern = 8'b00110000; 
    { 8'h3b, 4'hc }: pattern = 8'b00000000; 
    { 8'h3b, 4'hd }: pattern = 8'b00000000; 
    { 8'h3b, 4'he }: pattern = 8'b00000000; 
    { 8'h3b, 4'hf }: pattern = 8'b00000000; 

    { 8'h3c, 4'h0 }: pattern = 8'b00000000; 
    { 8'h3c, 4'h1 }: pattern = 8'b00000000; 
    { 8'h3c, 4'h2 }: pattern = 8'b00000000; 
    { 8'h3c, 4'h3 }: pattern = 8'b00000110; 
    { 8'h3c, 4'h4 }: pattern = 8'b00001100; 
    { 8'h3c, 4'h5 }: pattern = 8'b00011000; 
    { 8'h3c, 4'h6 }: pattern = 8'b00110000; 
    { 8'h3c, 4'h7 }: pattern = 8'b01100000; 
    { 8'h3c, 4'h8 }: pattern = 8'b00110000; 
    { 8'h3c, 4'h9 }: pattern = 8'b00011000; 
    { 8'h3c, 4'ha }: pattern = 8'b00001100; 
    { 8'h3c, 4'hb }: pattern = 8'b00000110; 
    { 8'h3c, 4'hc }: pattern = 8'b00000000; 
    { 8'h3c, 4'hd }: pattern = 8'b00000000; 
    { 8'h3c, 4'he }: pattern = 8'b00000000; 
    { 8'h3c, 4'hf }: pattern = 8'b00000000; 

    { 8'h3d, 4'h0 }: pattern = 8'b00000000; 
    { 8'h3d, 4'h1 }: pattern = 8'b00000000; 
    { 8'h3d, 4'h2 }: pattern = 8'b00000000; 
    { 8'h3d, 4'h3 }: pattern = 8'b00000000; 
    { 8'h3d, 4'h4 }: pattern = 8'b00000000; 
    { 8'h3d, 4'h5 }: pattern = 8'b01111110; 
    { 8'h3d, 4'h6 }: pattern = 8'b00000000; 
    { 8'h3d, 4'h7 }: pattern = 8'b00000000; 
    { 8'h3d, 4'h8 }: pattern = 8'b01111110; 
    { 8'h3d, 4'h9 }: pattern = 8'b00000000; 
    { 8'h3d, 4'ha }: pattern = 8'b00000000; 
    { 8'h3d, 4'hb }: pattern = 8'b00000000; 
    { 8'h3d, 4'hc }: pattern = 8'b00000000; 
    { 8'h3d, 4'hd }: pattern = 8'b00000000; 
    { 8'h3d, 4'he }: pattern = 8'b00000000; 
    { 8'h3d, 4'hf }: pattern = 8'b00000000; 

    { 8'h3e, 4'h0 }: pattern = 8'b00000000; 
    { 8'h3e, 4'h1 }: pattern = 8'b00000000; 
    { 8'h3e, 4'h2 }: pattern = 8'b00000000; 
    { 8'h3e, 4'h3 }: pattern = 8'b01100000; 
    { 8'h3e, 4'h4 }: pattern = 8'b00110000; 
    { 8'h3e, 4'h5 }: pattern = 8'b00011000; 
    { 8'h3e, 4'h6 }: pattern = 8'b00001100; 
    { 8'h3e, 4'h7 }: pattern = 8'b00000110; 
    { 8'h3e, 4'h8 }: pattern = 8'b00001100; 
    { 8'h3e, 4'h9 }: pattern = 8'b00011000; 
    { 8'h3e, 4'ha }: pattern = 8'b00110000; 
    { 8'h3e, 4'hb }: pattern = 8'b01100000; 
    { 8'h3e, 4'hc }: pattern = 8'b00000000; 
    { 8'h3e, 4'hd }: pattern = 8'b00000000; 
    { 8'h3e, 4'he }: pattern = 8'b00000000; 
    { 8'h3e, 4'hf }: pattern = 8'b00000000; 

    { 8'h3f, 4'h0 }: pattern = 8'b00000000; 
    { 8'h3f, 4'h1 }: pattern = 8'b00000000; 
    { 8'h3f, 4'h2 }: pattern = 8'b01111100; 
    { 8'h3f, 4'h3 }: pattern = 8'b11000110; 
    { 8'h3f, 4'h4 }: pattern = 8'b11000110; 
    { 8'h3f, 4'h5 }: pattern = 8'b00001100; 
    { 8'h3f, 4'h6 }: pattern = 8'b00011000; 
    { 8'h3f, 4'h7 }: pattern = 8'b00011000; 
    { 8'h3f, 4'h8 }: pattern = 8'b00011000; 
    { 8'h3f, 4'h9 }: pattern = 8'b00000000; 
    { 8'h3f, 4'ha }: pattern = 8'b00011000; 
    { 8'h3f, 4'hb }: pattern = 8'b00011000; 
    { 8'h3f, 4'hc }: pattern = 8'b00000000; 
    { 8'h3f, 4'hd }: pattern = 8'b00000000; 
    { 8'h3f, 4'he }: pattern = 8'b00000000; 
    { 8'h3f, 4'hf }: pattern = 8'b00000000; 

    { 8'h40, 4'h0 }: pattern = 8'b00000000; 
    { 8'h40, 4'h1 }: pattern = 8'b00000000; 
    { 8'h40, 4'h2 }: pattern = 8'b00000000; 
    { 8'h40, 4'h3 }: pattern = 8'b01111100; 
    { 8'h40, 4'h4 }: pattern = 8'b11000110; 
    { 8'h40, 4'h5 }: pattern = 8'b11000110; 
    { 8'h40, 4'h6 }: pattern = 8'b11011110; 
    { 8'h40, 4'h7 }: pattern = 8'b11011110; 
    { 8'h40, 4'h8 }: pattern = 8'b11011110; 
    { 8'h40, 4'h9 }: pattern = 8'b11011100; 
    { 8'h40, 4'ha }: pattern = 8'b11000000; 
    { 8'h40, 4'hb }: pattern = 8'b01111100; 
    { 8'h40, 4'hc }: pattern = 8'b00000000; 
    { 8'h40, 4'hd }: pattern = 8'b00000000; 
    { 8'h40, 4'he }: pattern = 8'b00000000; 
    { 8'h40, 4'hf }: pattern = 8'b00000000; 

    { 8'h41, 4'h0 }: pattern = 8'b00000000; 
    { 8'h41, 4'h1 }: pattern = 8'b00000000; 
    { 8'h41, 4'h2 }: pattern = 8'b00010000; 
    { 8'h41, 4'h3 }: pattern = 8'b00111000; 
    { 8'h41, 4'h4 }: pattern = 8'b01101100; 
    { 8'h41, 4'h5 }: pattern = 8'b11000110; 
    { 8'h41, 4'h6 }: pattern = 8'b11000110; 
    { 8'h41, 4'h7 }: pattern = 8'b11111110; 
    { 8'h41, 4'h8 }: pattern = 8'b11000110; 
    { 8'h41, 4'h9 }: pattern = 8'b11000110; 
    { 8'h41, 4'ha }: pattern = 8'b11000110; 
    { 8'h41, 4'hb }: pattern = 8'b11000110; 
    { 8'h41, 4'hc }: pattern = 8'b00000000; 
    { 8'h41, 4'hd }: pattern = 8'b00000000; 
    { 8'h41, 4'he }: pattern = 8'b00000000; 
    { 8'h41, 4'hf }: pattern = 8'b00000000; 

    { 8'h42, 4'h0 }: pattern = 8'b00000000; 
    { 8'h42, 4'h1 }: pattern = 8'b00000000; 
    { 8'h42, 4'h2 }: pattern = 8'b11111100; 
    { 8'h42, 4'h3 }: pattern = 8'b01100110; 
    { 8'h42, 4'h4 }: pattern = 8'b01100110; 
    { 8'h42, 4'h5 }: pattern = 8'b01100110; 
    { 8'h42, 4'h6 }: pattern = 8'b01111100; 
    { 8'h42, 4'h7 }: pattern = 8'b01100110; 
    { 8'h42, 4'h8 }: pattern = 8'b01100110; 
    { 8'h42, 4'h9 }: pattern = 8'b01100110; 
    { 8'h42, 4'ha }: pattern = 8'b01100110; 
    { 8'h42, 4'hb }: pattern = 8'b11111100; 
    { 8'h42, 4'hc }: pattern = 8'b00000000; 
    { 8'h42, 4'hd }: pattern = 8'b00000000; 
    { 8'h42, 4'he }: pattern = 8'b00000000; 
    { 8'h42, 4'hf }: pattern = 8'b00000000; 

    { 8'h43, 4'h0 }: pattern = 8'b00000000; 
    { 8'h43, 4'h1 }: pattern = 8'b00000000; 
    { 8'h43, 4'h2 }: pattern = 8'b00111100; 
    { 8'h43, 4'h3 }: pattern = 8'b01100110; 
    { 8'h43, 4'h4 }: pattern = 8'b11000010; 
    { 8'h43, 4'h5 }: pattern = 8'b11000000; 
    { 8'h43, 4'h6 }: pattern = 8'b11000000; 
    { 8'h43, 4'h7 }: pattern = 8'b11000000; 
    { 8'h43, 4'h8 }: pattern = 8'b11000000; 
    { 8'h43, 4'h9 }: pattern = 8'b11000010; 
    { 8'h43, 4'ha }: pattern = 8'b01100110; 
    { 8'h43, 4'hb }: pattern = 8'b00111100; 
    { 8'h43, 4'hc }: pattern = 8'b00000000; 
    { 8'h43, 4'hd }: pattern = 8'b00000000; 
    { 8'h43, 4'he }: pattern = 8'b00000000; 
    { 8'h43, 4'hf }: pattern = 8'b00000000; 

    { 8'h44, 4'h0 }: pattern = 8'b00000000; 
    { 8'h44, 4'h1 }: pattern = 8'b00000000; 
    { 8'h44, 4'h2 }: pattern = 8'b11111000; 
    { 8'h44, 4'h3 }: pattern = 8'b01101100; 
    { 8'h44, 4'h4 }: pattern = 8'b01100110; 
    { 8'h44, 4'h5 }: pattern = 8'b01100110; 
    { 8'h44, 4'h6 }: pattern = 8'b01100110; 
    { 8'h44, 4'h7 }: pattern = 8'b01100110; 
    { 8'h44, 4'h8 }: pattern = 8'b01100110; 
    { 8'h44, 4'h9 }: pattern = 8'b01100110; 
    { 8'h44, 4'ha }: pattern = 8'b01101100; 
    { 8'h44, 4'hb }: pattern = 8'b11111000; 
    { 8'h44, 4'hc }: pattern = 8'b00000000; 
    { 8'h44, 4'hd }: pattern = 8'b00000000; 
    { 8'h44, 4'he }: pattern = 8'b00000000; 
    { 8'h44, 4'hf }: pattern = 8'b00000000; 

    { 8'h45, 4'h0 }: pattern = 8'b00000000; 
    { 8'h45, 4'h1 }: pattern = 8'b00000000; 
    { 8'h45, 4'h2 }: pattern = 8'b11111110; 
    { 8'h45, 4'h3 }: pattern = 8'b01100110; 
    { 8'h45, 4'h4 }: pattern = 8'b01100010; 
    { 8'h45, 4'h5 }: pattern = 8'b01101000; 
    { 8'h45, 4'h6 }: pattern = 8'b01111000; 
    { 8'h45, 4'h7 }: pattern = 8'b01101000; 
    { 8'h45, 4'h8 }: pattern = 8'b01100000; 
    { 8'h45, 4'h9 }: pattern = 8'b01100010; 
    { 8'h45, 4'ha }: pattern = 8'b01100110; 
    { 8'h45, 4'hb }: pattern = 8'b11111110; 
    { 8'h45, 4'hc }: pattern = 8'b00000000; 
    { 8'h45, 4'hd }: pattern = 8'b00000000; 
    { 8'h45, 4'he }: pattern = 8'b00000000; 
    { 8'h45, 4'hf }: pattern = 8'b00000000; 

    { 8'h46, 4'h0 }: pattern = 8'b00000000; 
    { 8'h46, 4'h1 }: pattern = 8'b00000000; 
    { 8'h46, 4'h2 }: pattern = 8'b11111110; 
    { 8'h46, 4'h3 }: pattern = 8'b01100110; 
    { 8'h46, 4'h4 }: pattern = 8'b01100010; 
    { 8'h46, 4'h5 }: pattern = 8'b01101000; 
    { 8'h46, 4'h6 }: pattern = 8'b01111000; 
    { 8'h46, 4'h7 }: pattern = 8'b01101000; 
    { 8'h46, 4'h8 }: pattern = 8'b01100000; 
    { 8'h46, 4'h9 }: pattern = 8'b01100000; 
    { 8'h46, 4'ha }: pattern = 8'b01100000; 
    { 8'h46, 4'hb }: pattern = 8'b11110000; 
    { 8'h46, 4'hc }: pattern = 8'b00000000; 
    { 8'h46, 4'hd }: pattern = 8'b00000000; 
    { 8'h46, 4'he }: pattern = 8'b00000000; 
    { 8'h46, 4'hf }: pattern = 8'b00000000; 

    { 8'h47, 4'h0 }: pattern = 8'b00000000; 
    { 8'h47, 4'h1 }: pattern = 8'b00000000; 
    { 8'h47, 4'h2 }: pattern = 8'b00111100; 
    { 8'h47, 4'h3 }: pattern = 8'b01100110; 
    { 8'h47, 4'h4 }: pattern = 8'b11000010; 
    { 8'h47, 4'h5 }: pattern = 8'b11000000; 
    { 8'h47, 4'h6 }: pattern = 8'b11000000; 
    { 8'h47, 4'h7 }: pattern = 8'b11011110; 
    { 8'h47, 4'h8 }: pattern = 8'b11000110; 
    { 8'h47, 4'h9 }: pattern = 8'b11000110; 
    { 8'h47, 4'ha }: pattern = 8'b01100110; 
    { 8'h47, 4'hb }: pattern = 8'b00111010; 
    { 8'h47, 4'hc }: pattern = 8'b00000000; 
    { 8'h47, 4'hd }: pattern = 8'b00000000; 
    { 8'h47, 4'he }: pattern = 8'b00000000; 
    { 8'h47, 4'hf }: pattern = 8'b00000000; 

    { 8'h48, 4'h0 }: pattern = 8'b00000000; 
    { 8'h48, 4'h1 }: pattern = 8'b00000000; 
    { 8'h48, 4'h2 }: pattern = 8'b11000110; 
    { 8'h48, 4'h3 }: pattern = 8'b11000110; 
    { 8'h48, 4'h4 }: pattern = 8'b11000110; 
    { 8'h48, 4'h5 }: pattern = 8'b11000110; 
    { 8'h48, 4'h6 }: pattern = 8'b11111110; 
    { 8'h48, 4'h7 }: pattern = 8'b11000110; 
    { 8'h48, 4'h8 }: pattern = 8'b11000110; 
    { 8'h48, 4'h9 }: pattern = 8'b11000110; 
    { 8'h48, 4'ha }: pattern = 8'b11000110; 
    { 8'h48, 4'hb }: pattern = 8'b11000110; 
    { 8'h48, 4'hc }: pattern = 8'b00000000; 
    { 8'h48, 4'hd }: pattern = 8'b00000000; 
    { 8'h48, 4'he }: pattern = 8'b00000000; 
    { 8'h48, 4'hf }: pattern = 8'b00000000; 

    { 8'h49, 4'h0 }: pattern = 8'b00000000; 
    { 8'h49, 4'h1 }: pattern = 8'b00000000; 
    { 8'h49, 4'h2 }: pattern = 8'b00111100; 
    { 8'h49, 4'h3 }: pattern = 8'b00011000; 
    { 8'h49, 4'h4 }: pattern = 8'b00011000; 
    { 8'h49, 4'h5 }: pattern = 8'b00011000; 
    { 8'h49, 4'h6 }: pattern = 8'b00011000; 
    { 8'h49, 4'h7 }: pattern = 8'b00011000; 
    { 8'h49, 4'h8 }: pattern = 8'b00011000; 
    { 8'h49, 4'h9 }: pattern = 8'b00011000; 
    { 8'h49, 4'ha }: pattern = 8'b00011000; 
    { 8'h49, 4'hb }: pattern = 8'b00111100; 
    { 8'h49, 4'hc }: pattern = 8'b00000000; 
    { 8'h49, 4'hd }: pattern = 8'b00000000; 
    { 8'h49, 4'he }: pattern = 8'b00000000; 
    { 8'h49, 4'hf }: pattern = 8'b00000000; 

    { 8'h4a, 4'h0 }: pattern = 8'b00000000; 
    { 8'h4a, 4'h1 }: pattern = 8'b00000000; 
    { 8'h4a, 4'h2 }: pattern = 8'b00011110; 
    { 8'h4a, 4'h3 }: pattern = 8'b00001100; 
    { 8'h4a, 4'h4 }: pattern = 8'b00001100; 
    { 8'h4a, 4'h5 }: pattern = 8'b00001100; 
    { 8'h4a, 4'h6 }: pattern = 8'b00001100; 
    { 8'h4a, 4'h7 }: pattern = 8'b00001100; 
    { 8'h4a, 4'h8 }: pattern = 8'b11001100; 
    { 8'h4a, 4'h9 }: pattern = 8'b11001100; 
    { 8'h4a, 4'ha }: pattern = 8'b11001100; 
    { 8'h4a, 4'hb }: pattern = 8'b01111000; 
    { 8'h4a, 4'hc }: pattern = 8'b00000000; 
    { 8'h4a, 4'hd }: pattern = 8'b00000000; 
    { 8'h4a, 4'he }: pattern = 8'b00000000; 
    { 8'h4a, 4'hf }: pattern = 8'b00000000; 

    { 8'h4b, 4'h0 }: pattern = 8'b00000000; 
    { 8'h4b, 4'h1 }: pattern = 8'b00000000; 
    { 8'h4b, 4'h2 }: pattern = 8'b11100110; 
    { 8'h4b, 4'h3 }: pattern = 8'b01100110; 
    { 8'h4b, 4'h4 }: pattern = 8'b01100110; 
    { 8'h4b, 4'h5 }: pattern = 8'b01101100; 
    { 8'h4b, 4'h6 }: pattern = 8'b01111000; 
    { 8'h4b, 4'h7 }: pattern = 8'b01111000; 
    { 8'h4b, 4'h8 }: pattern = 8'b01101100; 
    { 8'h4b, 4'h9 }: pattern = 8'b01100110; 
    { 8'h4b, 4'ha }: pattern = 8'b01100110; 
    { 8'h4b, 4'hb }: pattern = 8'b11100110; 
    { 8'h4b, 4'hc }: pattern = 8'b00000000; 
    { 8'h4b, 4'hd }: pattern = 8'b00000000; 
    { 8'h4b, 4'he }: pattern = 8'b00000000; 
    { 8'h4b, 4'hf }: pattern = 8'b00000000; 

    { 8'h4c, 4'h0 }: pattern = 8'b00000000; 
    { 8'h4c, 4'h1 }: pattern = 8'b00000000; 
    { 8'h4c, 4'h2 }: pattern = 8'b11110000; 
    { 8'h4c, 4'h3 }: pattern = 8'b01100000; 
    { 8'h4c, 4'h4 }: pattern = 8'b01100000; 
    { 8'h4c, 4'h5 }: pattern = 8'b01100000; 
    { 8'h4c, 4'h6 }: pattern = 8'b01100000; 
    { 8'h4c, 4'h7 }: pattern = 8'b01100000; 
    { 8'h4c, 4'h8 }: pattern = 8'b01100000; 
    { 8'h4c, 4'h9 }: pattern = 8'b01100010; 
    { 8'h4c, 4'ha }: pattern = 8'b01100110; 
    { 8'h4c, 4'hb }: pattern = 8'b11111110; 
    { 8'h4c, 4'hc }: pattern = 8'b00000000; 
    { 8'h4c, 4'hd }: pattern = 8'b00000000; 
    { 8'h4c, 4'he }: pattern = 8'b00000000; 
    { 8'h4c, 4'hf }: pattern = 8'b00000000; 

    { 8'h4d, 4'h0 }: pattern = 8'b00000000; 
    { 8'h4d, 4'h1 }: pattern = 8'b00000000; 
    { 8'h4d, 4'h2 }: pattern = 8'b11000110; 
    { 8'h4d, 4'h3 }: pattern = 8'b11101110; 
    { 8'h4d, 4'h4 }: pattern = 8'b11111110; 
    { 8'h4d, 4'h5 }: pattern = 8'b11111110; 
    { 8'h4d, 4'h6 }: pattern = 8'b11010110; 
    { 8'h4d, 4'h7 }: pattern = 8'b11000110; 
    { 8'h4d, 4'h8 }: pattern = 8'b11000110; 
    { 8'h4d, 4'h9 }: pattern = 8'b11000110; 
    { 8'h4d, 4'ha }: pattern = 8'b11000110; 
    { 8'h4d, 4'hb }: pattern = 8'b11000110; 
    { 8'h4d, 4'hc }: pattern = 8'b00000000; 
    { 8'h4d, 4'hd }: pattern = 8'b00000000; 
    { 8'h4d, 4'he }: pattern = 8'b00000000; 
    { 8'h4d, 4'hf }: pattern = 8'b00000000; 

    { 8'h4e, 4'h0 }: pattern = 8'b00000000; 
    { 8'h4e, 4'h1 }: pattern = 8'b00000000; 
    { 8'h4e, 4'h2 }: pattern = 8'b11000110; 
    { 8'h4e, 4'h3 }: pattern = 8'b11100110; 
    { 8'h4e, 4'h4 }: pattern = 8'b11110110; 
    { 8'h4e, 4'h5 }: pattern = 8'b11111110; 
    { 8'h4e, 4'h6 }: pattern = 8'b11011110; 
    { 8'h4e, 4'h7 }: pattern = 8'b11001110; 
    { 8'h4e, 4'h8 }: pattern = 8'b11000110; 
    { 8'h4e, 4'h9 }: pattern = 8'b11000110; 
    { 8'h4e, 4'ha }: pattern = 8'b11000110; 
    { 8'h4e, 4'hb }: pattern = 8'b11000110; 
    { 8'h4e, 4'hc }: pattern = 8'b00000000; 
    { 8'h4e, 4'hd }: pattern = 8'b00000000; 
    { 8'h4e, 4'he }: pattern = 8'b00000000; 
    { 8'h4e, 4'hf }: pattern = 8'b00000000; 

    { 8'h4f, 4'h0 }: pattern = 8'b00000000; 
    { 8'h4f, 4'h1 }: pattern = 8'b00000000; 
    { 8'h4f, 4'h2 }: pattern = 8'b01111100; 
    { 8'h4f, 4'h3 }: pattern = 8'b11000110; 
    { 8'h4f, 4'h4 }: pattern = 8'b11000110; 
    { 8'h4f, 4'h5 }: pattern = 8'b11000110; 
    { 8'h4f, 4'h6 }: pattern = 8'b11000110; 
    { 8'h4f, 4'h7 }: pattern = 8'b11000110; 
    { 8'h4f, 4'h8 }: pattern = 8'b11000110; 
    { 8'h4f, 4'h9 }: pattern = 8'b11000110; 
    { 8'h4f, 4'ha }: pattern = 8'b11000110; 
    { 8'h4f, 4'hb }: pattern = 8'b01111100; 
    { 8'h4f, 4'hc }: pattern = 8'b00000000; 
    { 8'h4f, 4'hd }: pattern = 8'b00000000; 
    { 8'h4f, 4'he }: pattern = 8'b00000000; 
    { 8'h4f, 4'hf }: pattern = 8'b00000000; 

    { 8'h50, 4'h0 }: pattern = 8'b00000000; 
    { 8'h50, 4'h1 }: pattern = 8'b00000000; 
    { 8'h50, 4'h2 }: pattern = 8'b11111100; 
    { 8'h50, 4'h3 }: pattern = 8'b01100110; 
    { 8'h50, 4'h4 }: pattern = 8'b01100110; 
    { 8'h50, 4'h5 }: pattern = 8'b01100110; 
    { 8'h50, 4'h6 }: pattern = 8'b01111100; 
    { 8'h50, 4'h7 }: pattern = 8'b01100000; 
    { 8'h50, 4'h8 }: pattern = 8'b01100000; 
    { 8'h50, 4'h9 }: pattern = 8'b01100000; 
    { 8'h50, 4'ha }: pattern = 8'b01100000; 
    { 8'h50, 4'hb }: pattern = 8'b11110000; 
    { 8'h50, 4'hc }: pattern = 8'b00000000; 
    { 8'h50, 4'hd }: pattern = 8'b00000000; 
    { 8'h50, 4'he }: pattern = 8'b00000000; 
    { 8'h50, 4'hf }: pattern = 8'b00000000; 

    { 8'h51, 4'h0 }: pattern = 8'b00000000; 
    { 8'h51, 4'h1 }: pattern = 8'b00000000; 
    { 8'h51, 4'h2 }: pattern = 8'b01111100; 
    { 8'h51, 4'h3 }: pattern = 8'b11000110; 
    { 8'h51, 4'h4 }: pattern = 8'b11000110; 
    { 8'h51, 4'h5 }: pattern = 8'b11000110; 
    { 8'h51, 4'h6 }: pattern = 8'b11000110; 
    { 8'h51, 4'h7 }: pattern = 8'b11000110; 
    { 8'h51, 4'h8 }: pattern = 8'b11000110; 
    { 8'h51, 4'h9 }: pattern = 8'b11010110; 
    { 8'h51, 4'ha }: pattern = 8'b11011110; 
    { 8'h51, 4'hb }: pattern = 8'b01111100; 
    { 8'h51, 4'hc }: pattern = 8'b00001100; 
    { 8'h51, 4'hd }: pattern = 8'b00001110; 
    { 8'h51, 4'he }: pattern = 8'b00000000; 
    { 8'h51, 4'hf }: pattern = 8'b00000000; 

    { 8'h52, 4'h0 }: pattern = 8'b00000000; 
    { 8'h52, 4'h1 }: pattern = 8'b00000000; 
    { 8'h52, 4'h2 }: pattern = 8'b11111100; 
    { 8'h52, 4'h3 }: pattern = 8'b01100110; 
    { 8'h52, 4'h4 }: pattern = 8'b01100110; 
    { 8'h52, 4'h5 }: pattern = 8'b01100110; 
    { 8'h52, 4'h6 }: pattern = 8'b01111100; 
    { 8'h52, 4'h7 }: pattern = 8'b01101100; 
    { 8'h52, 4'h8 }: pattern = 8'b01100110; 
    { 8'h52, 4'h9 }: pattern = 8'b01100110; 
    { 8'h52, 4'ha }: pattern = 8'b01100110; 
    { 8'h52, 4'hb }: pattern = 8'b11100110; 
    { 8'h52, 4'hc }: pattern = 8'b00000000; 
    { 8'h52, 4'hd }: pattern = 8'b00000000; 
    { 8'h52, 4'he }: pattern = 8'b00000000; 
    { 8'h52, 4'hf }: pattern = 8'b00000000; 

    { 8'h53, 4'h0 }: pattern = 8'b00000000; 
    { 8'h53, 4'h1 }: pattern = 8'b00000000; 
    { 8'h53, 4'h2 }: pattern = 8'b01111100; 
    { 8'h53, 4'h3 }: pattern = 8'b11000110; 
    { 8'h53, 4'h4 }: pattern = 8'b11000110; 
    { 8'h53, 4'h5 }: pattern = 8'b01100000; 
    { 8'h53, 4'h6 }: pattern = 8'b00111000; 
    { 8'h53, 4'h7 }: pattern = 8'b00001100; 
    { 8'h53, 4'h8 }: pattern = 8'b00000110; 
    { 8'h53, 4'h9 }: pattern = 8'b11000110; 
    { 8'h53, 4'ha }: pattern = 8'b11000110; 
    { 8'h53, 4'hb }: pattern = 8'b01111100; 
    { 8'h53, 4'hc }: pattern = 8'b00000000; 
    { 8'h53, 4'hd }: pattern = 8'b00000000; 
    { 8'h53, 4'he }: pattern = 8'b00000000; 
    { 8'h53, 4'hf }: pattern = 8'b00000000; 

    { 8'h54, 4'h0 }: pattern = 8'b00000000; 
    { 8'h54, 4'h1 }: pattern = 8'b00000000; 
    { 8'h54, 4'h2 }: pattern = 8'b01111110; 
    { 8'h54, 4'h3 }: pattern = 8'b01111110; 
    { 8'h54, 4'h4 }: pattern = 8'b01011010; 
    { 8'h54, 4'h5 }: pattern = 8'b00011000; 
    { 8'h54, 4'h6 }: pattern = 8'b00011000; 
    { 8'h54, 4'h7 }: pattern = 8'b00011000; 
    { 8'h54, 4'h8 }: pattern = 8'b00011000; 
    { 8'h54, 4'h9 }: pattern = 8'b00011000; 
    { 8'h54, 4'ha }: pattern = 8'b00011000; 
    { 8'h54, 4'hb }: pattern = 8'b00111100; 
    { 8'h54, 4'hc }: pattern = 8'b00000000; 
    { 8'h54, 4'hd }: pattern = 8'b00000000; 
    { 8'h54, 4'he }: pattern = 8'b00000000; 
    { 8'h54, 4'hf }: pattern = 8'b00000000; 

    { 8'h55, 4'h0 }: pattern = 8'b00000000; 
    { 8'h55, 4'h1 }: pattern = 8'b00000000; 
    { 8'h55, 4'h2 }: pattern = 8'b11000110; 
    { 8'h55, 4'h3 }: pattern = 8'b11000110; 
    { 8'h55, 4'h4 }: pattern = 8'b11000110; 
    { 8'h55, 4'h5 }: pattern = 8'b11000110; 
    { 8'h55, 4'h6 }: pattern = 8'b11000110; 
    { 8'h55, 4'h7 }: pattern = 8'b11000110; 
    { 8'h55, 4'h8 }: pattern = 8'b11000110; 
    { 8'h55, 4'h9 }: pattern = 8'b11000110; 
    { 8'h55, 4'ha }: pattern = 8'b11000110; 
    { 8'h55, 4'hb }: pattern = 8'b01111100; 
    { 8'h55, 4'hc }: pattern = 8'b00000000; 
    { 8'h55, 4'hd }: pattern = 8'b00000000; 
    { 8'h55, 4'he }: pattern = 8'b00000000; 
    { 8'h55, 4'hf }: pattern = 8'b00000000; 

    { 8'h56, 4'h0 }: pattern = 8'b00000000; 
    { 8'h56, 4'h1 }: pattern = 8'b00000000; 
    { 8'h56, 4'h2 }: pattern = 8'b11000110; 
    { 8'h56, 4'h3 }: pattern = 8'b11000110; 
    { 8'h56, 4'h4 }: pattern = 8'b11000110; 
    { 8'h56, 4'h5 }: pattern = 8'b11000110; 
    { 8'h56, 4'h6 }: pattern = 8'b11000110; 
    { 8'h56, 4'h7 }: pattern = 8'b11000110; 
    { 8'h56, 4'h8 }: pattern = 8'b11000110; 
    { 8'h56, 4'h9 }: pattern = 8'b01101100; 
    { 8'h56, 4'ha }: pattern = 8'b00111000; 
    { 8'h56, 4'hb }: pattern = 8'b00010000; 
    { 8'h56, 4'hc }: pattern = 8'b00000000; 
    { 8'h56, 4'hd }: pattern = 8'b00000000; 
    { 8'h56, 4'he }: pattern = 8'b00000000; 
    { 8'h56, 4'hf }: pattern = 8'b00000000; 

    { 8'h57, 4'h0 }: pattern = 8'b00000000; 
    { 8'h57, 4'h1 }: pattern = 8'b00000000; 
    { 8'h57, 4'h2 }: pattern = 8'b11000110; 
    { 8'h57, 4'h3 }: pattern = 8'b11000110; 
    { 8'h57, 4'h4 }: pattern = 8'b11000110; 
    { 8'h57, 4'h5 }: pattern = 8'b11000110; 
    { 8'h57, 4'h6 }: pattern = 8'b11010110; 
    { 8'h57, 4'h7 }: pattern = 8'b11010110; 
    { 8'h57, 4'h8 }: pattern = 8'b11010110; 
    { 8'h57, 4'h9 }: pattern = 8'b11111110; 
    { 8'h57, 4'ha }: pattern = 8'b11101110; 
    { 8'h57, 4'hb }: pattern = 8'b01101100; 
    { 8'h57, 4'hc }: pattern = 8'b00000000; 
    { 8'h57, 4'hd }: pattern = 8'b00000000; 
    { 8'h57, 4'he }: pattern = 8'b00000000; 
    { 8'h57, 4'hf }: pattern = 8'b00000000; 

    { 8'h58, 4'h0 }: pattern = 8'b00000000; 
    { 8'h58, 4'h1 }: pattern = 8'b00000000; 
    { 8'h58, 4'h2 }: pattern = 8'b11000110; 
    { 8'h58, 4'h3 }: pattern = 8'b11000110; 
    { 8'h58, 4'h4 }: pattern = 8'b01101100; 
    { 8'h58, 4'h5 }: pattern = 8'b01111100; 
    { 8'h58, 4'h6 }: pattern = 8'b00111000; 
    { 8'h58, 4'h7 }: pattern = 8'b00111000; 
    { 8'h58, 4'h8 }: pattern = 8'b01111100; 
    { 8'h58, 4'h9 }: pattern = 8'b01101100; 
    { 8'h58, 4'ha }: pattern = 8'b11000110; 
    { 8'h58, 4'hb }: pattern = 8'b11000110; 
    { 8'h58, 4'hc }: pattern = 8'b00000000; 
    { 8'h58, 4'hd }: pattern = 8'b00000000; 
    { 8'h58, 4'he }: pattern = 8'b00000000; 
    { 8'h58, 4'hf }: pattern = 8'b00000000; 

    { 8'h59, 4'h0 }: pattern = 8'b00000000; 
    { 8'h59, 4'h1 }: pattern = 8'b00000000; 
    { 8'h59, 4'h2 }: pattern = 8'b01100110; 
    { 8'h59, 4'h3 }: pattern = 8'b01100110; 
    { 8'h59, 4'h4 }: pattern = 8'b01100110; 
    { 8'h59, 4'h5 }: pattern = 8'b01100110; 
    { 8'h59, 4'h6 }: pattern = 8'b00111100; 
    { 8'h59, 4'h7 }: pattern = 8'b00011000; 
    { 8'h59, 4'h8 }: pattern = 8'b00011000; 
    { 8'h59, 4'h9 }: pattern = 8'b00011000; 
    { 8'h59, 4'ha }: pattern = 8'b00011000; 
    { 8'h59, 4'hb }: pattern = 8'b00111100; 
    { 8'h59, 4'hc }: pattern = 8'b00000000; 
    { 8'h59, 4'hd }: pattern = 8'b00000000; 
    { 8'h59, 4'he }: pattern = 8'b00000000; 
    { 8'h59, 4'hf }: pattern = 8'b00000000; 

    { 8'h5a, 4'h0 }: pattern = 8'b00000000; 
    { 8'h5a, 4'h1 }: pattern = 8'b00000000; 
    { 8'h5a, 4'h2 }: pattern = 8'b11111110; 
    { 8'h5a, 4'h3 }: pattern = 8'b11000110; 
    { 8'h5a, 4'h4 }: pattern = 8'b10000110; 
    { 8'h5a, 4'h5 }: pattern = 8'b00001100; 
    { 8'h5a, 4'h6 }: pattern = 8'b00011000; 
    { 8'h5a, 4'h7 }: pattern = 8'b00110000; 
    { 8'h5a, 4'h8 }: pattern = 8'b01100000; 
    { 8'h5a, 4'h9 }: pattern = 8'b11000010; 
    { 8'h5a, 4'ha }: pattern = 8'b11000110; 
    { 8'h5a, 4'hb }: pattern = 8'b11111110; 
    { 8'h5a, 4'hc }: pattern = 8'b00000000; 
    { 8'h5a, 4'hd }: pattern = 8'b00000000; 
    { 8'h5a, 4'he }: pattern = 8'b00000000; 
    { 8'h5a, 4'hf }: pattern = 8'b00000000; 

    { 8'h5b, 4'h0 }: pattern = 8'b00000000; 
    { 8'h5b, 4'h1 }: pattern = 8'b00000000; 
    { 8'h5b, 4'h2 }: pattern = 8'b00111100; 
    { 8'h5b, 4'h3 }: pattern = 8'b00110000; 
    { 8'h5b, 4'h4 }: pattern = 8'b00110000; 
    { 8'h5b, 4'h5 }: pattern = 8'b00110000; 
    { 8'h5b, 4'h6 }: pattern = 8'b00110000; 
    { 8'h5b, 4'h7 }: pattern = 8'b00110000; 
    { 8'h5b, 4'h8 }: pattern = 8'b00110000; 
    { 8'h5b, 4'h9 }: pattern = 8'b00110000; 
    { 8'h5b, 4'ha }: pattern = 8'b00110000; 
    { 8'h5b, 4'hb }: pattern = 8'b00111100; 
    { 8'h5b, 4'hc }: pattern = 8'b00000000; 
    { 8'h5b, 4'hd }: pattern = 8'b00000000; 
    { 8'h5b, 4'he }: pattern = 8'b00000000; 
    { 8'h5b, 4'hf }: pattern = 8'b00000000; 

    { 8'h5c, 4'h0 }: pattern = 8'b00000000; 
    { 8'h5c, 4'h1 }: pattern = 8'b00000000; 
    { 8'h5c, 4'h2 }: pattern = 8'b00000000; 
    { 8'h5c, 4'h3 }: pattern = 8'b10000000; 
    { 8'h5c, 4'h4 }: pattern = 8'b11000000; 
    { 8'h5c, 4'h5 }: pattern = 8'b11100000; 
    { 8'h5c, 4'h6 }: pattern = 8'b01110000; 
    { 8'h5c, 4'h7 }: pattern = 8'b00111000; 
    { 8'h5c, 4'h8 }: pattern = 8'b00011100; 
    { 8'h5c, 4'h9 }: pattern = 8'b00001110; 
    { 8'h5c, 4'ha }: pattern = 8'b00000110; 
    { 8'h5c, 4'hb }: pattern = 8'b00000010; 
    { 8'h5c, 4'hc }: pattern = 8'b00000000; 
    { 8'h5c, 4'hd }: pattern = 8'b00000000; 
    { 8'h5c, 4'he }: pattern = 8'b00000000; 
    { 8'h5c, 4'hf }: pattern = 8'b00000000; 

    { 8'h5d, 4'h0 }: pattern = 8'b00000000; 
    { 8'h5d, 4'h1 }: pattern = 8'b00000000; 
    { 8'h5d, 4'h2 }: pattern = 8'b00111100; 
    { 8'h5d, 4'h3 }: pattern = 8'b00001100; 
    { 8'h5d, 4'h4 }: pattern = 8'b00001100; 
    { 8'h5d, 4'h5 }: pattern = 8'b00001100; 
    { 8'h5d, 4'h6 }: pattern = 8'b00001100; 
    { 8'h5d, 4'h7 }: pattern = 8'b00001100; 
    { 8'h5d, 4'h8 }: pattern = 8'b00001100; 
    { 8'h5d, 4'h9 }: pattern = 8'b00001100; 
    { 8'h5d, 4'ha }: pattern = 8'b00001100; 
    { 8'h5d, 4'hb }: pattern = 8'b00111100; 
    { 8'h5d, 4'hc }: pattern = 8'b00000000; 
    { 8'h5d, 4'hd }: pattern = 8'b00000000; 
    { 8'h5d, 4'he }: pattern = 8'b00000000; 
    { 8'h5d, 4'hf }: pattern = 8'b00000000; 

    { 8'h5e, 4'h0 }: pattern = 8'b00010000; 
    { 8'h5e, 4'h1 }: pattern = 8'b00111000; 
    { 8'h5e, 4'h2 }: pattern = 8'b01101100; 
    { 8'h5e, 4'h3 }: pattern = 8'b11000110; 
    { 8'h5e, 4'h4 }: pattern = 8'b00000000; 
    { 8'h5e, 4'h5 }: pattern = 8'b00000000; 
    { 8'h5e, 4'h6 }: pattern = 8'b00000000; 
    { 8'h5e, 4'h7 }: pattern = 8'b00000000; 
    { 8'h5e, 4'h8 }: pattern = 8'b00000000; 
    { 8'h5e, 4'h9 }: pattern = 8'b00000000; 
    { 8'h5e, 4'ha }: pattern = 8'b00000000; 
    { 8'h5e, 4'hb }: pattern = 8'b00000000; 
    { 8'h5e, 4'hc }: pattern = 8'b00000000; 
    { 8'h5e, 4'hd }: pattern = 8'b00000000; 
    { 8'h5e, 4'he }: pattern = 8'b00000000; 
    { 8'h5e, 4'hf }: pattern = 8'b00000000; 

    { 8'h5f, 4'h0 }: pattern = 8'b00000000; 
    { 8'h5f, 4'h1 }: pattern = 8'b00000000; 
    { 8'h5f, 4'h2 }: pattern = 8'b00000000; 
    { 8'h5f, 4'h3 }: pattern = 8'b00000000; 
    { 8'h5f, 4'h4 }: pattern = 8'b00000000; 
    { 8'h5f, 4'h5 }: pattern = 8'b00000000; 
    { 8'h5f, 4'h6 }: pattern = 8'b00000000; 
    { 8'h5f, 4'h7 }: pattern = 8'b00000000; 
    { 8'h5f, 4'h8 }: pattern = 8'b00000000; 
    { 8'h5f, 4'h9 }: pattern = 8'b00000000; 
    { 8'h5f, 4'ha }: pattern = 8'b00000000; 
    { 8'h5f, 4'hb }: pattern = 8'b00000000; 
    { 8'h5f, 4'hc }: pattern = 8'b00000000; 
    { 8'h5f, 4'hd }: pattern = 8'b11111111; 
    { 8'h5f, 4'he }: pattern = 8'b00000000; 
    { 8'h5f, 4'hf }: pattern = 8'b00000000; 

    { 8'h60, 4'h0 }: pattern = 8'b00110000; 
    { 8'h60, 4'h1 }: pattern = 8'b00110000; 
    { 8'h60, 4'h2 }: pattern = 8'b00011000; 
    { 8'h60, 4'h3 }: pattern = 8'b00000000; 
    { 8'h60, 4'h4 }: pattern = 8'b00000000; 
    { 8'h60, 4'h5 }: pattern = 8'b00000000; 
    { 8'h60, 4'h6 }: pattern = 8'b00000000; 
    { 8'h60, 4'h7 }: pattern = 8'b00000000; 
    { 8'h60, 4'h8 }: pattern = 8'b00000000; 
    { 8'h60, 4'h9 }: pattern = 8'b00000000; 
    { 8'h60, 4'ha }: pattern = 8'b00000000; 
    { 8'h60, 4'hb }: pattern = 8'b00000000; 
    { 8'h60, 4'hc }: pattern = 8'b00000000; 
    { 8'h60, 4'hd }: pattern = 8'b00000000; 
    { 8'h60, 4'he }: pattern = 8'b00000000; 
    { 8'h60, 4'hf }: pattern = 8'b00000000; 

    { 8'h61, 4'h0 }: pattern = 8'b00000000; 
    { 8'h61, 4'h1 }: pattern = 8'b00000000; 
    { 8'h61, 4'h2 }: pattern = 8'b00000000; 
    { 8'h61, 4'h3 }: pattern = 8'b00000000; 
    { 8'h61, 4'h4 }: pattern = 8'b00000000; 
    { 8'h61, 4'h5 }: pattern = 8'b01111000; 
    { 8'h61, 4'h6 }: pattern = 8'b00001100; 
    { 8'h61, 4'h7 }: pattern = 8'b01111100; 
    { 8'h61, 4'h8 }: pattern = 8'b11001100; 
    { 8'h61, 4'h9 }: pattern = 8'b11001100; 
    { 8'h61, 4'ha }: pattern = 8'b11001100; 
    { 8'h61, 4'hb }: pattern = 8'b01110110; 
    { 8'h61, 4'hc }: pattern = 8'b00000000; 
    { 8'h61, 4'hd }: pattern = 8'b00000000; 
    { 8'h61, 4'he }: pattern = 8'b00000000; 
    { 8'h61, 4'hf }: pattern = 8'b00000000; 

    { 8'h62, 4'h0 }: pattern = 8'b00000000; 
    { 8'h62, 4'h1 }: pattern = 8'b00000000; 
    { 8'h62, 4'h2 }: pattern = 8'b11100000; 
    { 8'h62, 4'h3 }: pattern = 8'b01100000; 
    { 8'h62, 4'h4 }: pattern = 8'b01100000; 
    { 8'h62, 4'h5 }: pattern = 8'b01111000; 
    { 8'h62, 4'h6 }: pattern = 8'b01101100; 
    { 8'h62, 4'h7 }: pattern = 8'b01100110; 
    { 8'h62, 4'h8 }: pattern = 8'b01100110; 
    { 8'h62, 4'h9 }: pattern = 8'b01100110; 
    { 8'h62, 4'ha }: pattern = 8'b01100110; 
    { 8'h62, 4'hb }: pattern = 8'b01111100; 
    { 8'h62, 4'hc }: pattern = 8'b00000000; 
    { 8'h62, 4'hd }: pattern = 8'b00000000; 
    { 8'h62, 4'he }: pattern = 8'b00000000; 
    { 8'h62, 4'hf }: pattern = 8'b00000000; 

    { 8'h63, 4'h0 }: pattern = 8'b00000000; 
    { 8'h63, 4'h1 }: pattern = 8'b00000000; 
    { 8'h63, 4'h2 }: pattern = 8'b00000000; 
    { 8'h63, 4'h3 }: pattern = 8'b00000000; 
    { 8'h63, 4'h4 }: pattern = 8'b00000000; 
    { 8'h63, 4'h5 }: pattern = 8'b01111100; 
    { 8'h63, 4'h6 }: pattern = 8'b11000110; 
    { 8'h63, 4'h7 }: pattern = 8'b11000000; 
    { 8'h63, 4'h8 }: pattern = 8'b11000000; 
    { 8'h63, 4'h9 }: pattern = 8'b11000000; 
    { 8'h63, 4'ha }: pattern = 8'b11000110; 
    { 8'h63, 4'hb }: pattern = 8'b01111100; 
    { 8'h63, 4'hc }: pattern = 8'b00000000; 
    { 8'h63, 4'hd }: pattern = 8'b00000000; 
    { 8'h63, 4'he }: pattern = 8'b00000000; 
    { 8'h63, 4'hf }: pattern = 8'b00000000; 

    { 8'h64, 4'h0 }: pattern = 8'b00000000; 
    { 8'h64, 4'h1 }: pattern = 8'b00000000; 
    { 8'h64, 4'h2 }: pattern = 8'b00011100; 
    { 8'h64, 4'h3 }: pattern = 8'b00001100; 
    { 8'h64, 4'h4 }: pattern = 8'b00001100; 
    { 8'h64, 4'h5 }: pattern = 8'b00111100; 
    { 8'h64, 4'h6 }: pattern = 8'b01101100; 
    { 8'h64, 4'h7 }: pattern = 8'b11001100; 
    { 8'h64, 4'h8 }: pattern = 8'b11001100; 
    { 8'h64, 4'h9 }: pattern = 8'b11001100; 
    { 8'h64, 4'ha }: pattern = 8'b11001100; 
    { 8'h64, 4'hb }: pattern = 8'b01110110; 
    { 8'h64, 4'hc }: pattern = 8'b00000000; 
    { 8'h64, 4'hd }: pattern = 8'b00000000; 
    { 8'h64, 4'he }: pattern = 8'b00000000; 
    { 8'h64, 4'hf }: pattern = 8'b00000000; 

    { 8'h65, 4'h0 }: pattern = 8'b00000000; 
    { 8'h65, 4'h1 }: pattern = 8'b00000000; 
    { 8'h65, 4'h2 }: pattern = 8'b00000000; 
    { 8'h65, 4'h3 }: pattern = 8'b00000000; 
    { 8'h65, 4'h4 }: pattern = 8'b00000000; 
    { 8'h65, 4'h5 }: pattern = 8'b01111100; 
    { 8'h65, 4'h6 }: pattern = 8'b11000110; 
    { 8'h65, 4'h7 }: pattern = 8'b11111110; 
    { 8'h65, 4'h8 }: pattern = 8'b11000000; 
    { 8'h65, 4'h9 }: pattern = 8'b11000000; 
    { 8'h65, 4'ha }: pattern = 8'b11000110; 
    { 8'h65, 4'hb }: pattern = 8'b01111100; 
    { 8'h65, 4'hc }: pattern = 8'b00000000; 
    { 8'h65, 4'hd }: pattern = 8'b00000000; 
    { 8'h65, 4'he }: pattern = 8'b00000000; 
    { 8'h65, 4'hf }: pattern = 8'b00000000; 

    { 8'h66, 4'h0 }: pattern = 8'b00000000; 
    { 8'h66, 4'h1 }: pattern = 8'b00000000; 
    { 8'h66, 4'h2 }: pattern = 8'b00111000; 
    { 8'h66, 4'h3 }: pattern = 8'b01101100; 
    { 8'h66, 4'h4 }: pattern = 8'b01100100; 
    { 8'h66, 4'h5 }: pattern = 8'b01100000; 
    { 8'h66, 4'h6 }: pattern = 8'b11110000; 
    { 8'h66, 4'h7 }: pattern = 8'b01100000; 
    { 8'h66, 4'h8 }: pattern = 8'b01100000; 
    { 8'h66, 4'h9 }: pattern = 8'b01100000; 
    { 8'h66, 4'ha }: pattern = 8'b01100000; 
    { 8'h66, 4'hb }: pattern = 8'b11110000; 
    { 8'h66, 4'hc }: pattern = 8'b00000000; 
    { 8'h66, 4'hd }: pattern = 8'b00000000; 
    { 8'h66, 4'he }: pattern = 8'b00000000; 
    { 8'h66, 4'hf }: pattern = 8'b00000000; 

    { 8'h67, 4'h0 }: pattern = 8'b00000000; 
    { 8'h67, 4'h1 }: pattern = 8'b00000000; 
    { 8'h67, 4'h2 }: pattern = 8'b00000000; 
    { 8'h67, 4'h3 }: pattern = 8'b00000000; 
    { 8'h67, 4'h4 }: pattern = 8'b00000000; 
    { 8'h67, 4'h5 }: pattern = 8'b01110110; 
    { 8'h67, 4'h6 }: pattern = 8'b11001100; 
    { 8'h67, 4'h7 }: pattern = 8'b11001100; 
    { 8'h67, 4'h8 }: pattern = 8'b11001100; 
    { 8'h67, 4'h9 }: pattern = 8'b11001100; 
    { 8'h67, 4'ha }: pattern = 8'b11001100; 
    { 8'h67, 4'hb }: pattern = 8'b01111100; 
    { 8'h67, 4'hc }: pattern = 8'b00001100; 
    { 8'h67, 4'hd }: pattern = 8'b11001100; 
    { 8'h67, 4'he }: pattern = 8'b01111000; 
    { 8'h67, 4'hf }: pattern = 8'b00000000; 

    { 8'h68, 4'h0 }: pattern = 8'b00000000; 
    { 8'h68, 4'h1 }: pattern = 8'b00000000; 
    { 8'h68, 4'h2 }: pattern = 8'b11100000; 
    { 8'h68, 4'h3 }: pattern = 8'b01100000; 
    { 8'h68, 4'h4 }: pattern = 8'b01100000; 
    { 8'h68, 4'h5 }: pattern = 8'b01101100; 
    { 8'h68, 4'h6 }: pattern = 8'b01110110; 
    { 8'h68, 4'h7 }: pattern = 8'b01100110; 
    { 8'h68, 4'h8 }: pattern = 8'b01100110; 
    { 8'h68, 4'h9 }: pattern = 8'b01100110; 
    { 8'h68, 4'ha }: pattern = 8'b01100110; 
    { 8'h68, 4'hb }: pattern = 8'b11100110; 
    { 8'h68, 4'hc }: pattern = 8'b00000000; 
    { 8'h68, 4'hd }: pattern = 8'b00000000; 
    { 8'h68, 4'he }: pattern = 8'b00000000; 
    { 8'h68, 4'hf }: pattern = 8'b00000000; 

    { 8'h69, 4'h0 }: pattern = 8'b00000000; 
    { 8'h69, 4'h1 }: pattern = 8'b00000000; 
    { 8'h69, 4'h2 }: pattern = 8'b00011000; 
    { 8'h69, 4'h3 }: pattern = 8'b00011000; 
    { 8'h69, 4'h4 }: pattern = 8'b00000000; 
    { 8'h69, 4'h5 }: pattern = 8'b00111000; 
    { 8'h69, 4'h6 }: pattern = 8'b00011000; 
    { 8'h69, 4'h7 }: pattern = 8'b00011000; 
    { 8'h69, 4'h8 }: pattern = 8'b00011000; 
    { 8'h69, 4'h9 }: pattern = 8'b00011000; 
    { 8'h69, 4'ha }: pattern = 8'b00011000; 
    { 8'h69, 4'hb }: pattern = 8'b00111100; 
    { 8'h69, 4'hc }: pattern = 8'b00000000; 
    { 8'h69, 4'hd }: pattern = 8'b00000000; 
    { 8'h69, 4'he }: pattern = 8'b00000000; 
    { 8'h69, 4'hf }: pattern = 8'b00000000; 

    { 8'h6a, 4'h0 }: pattern = 8'b00000000; 
    { 8'h6a, 4'h1 }: pattern = 8'b00000000; 
    { 8'h6a, 4'h2 }: pattern = 8'b00000110; 
    { 8'h6a, 4'h3 }: pattern = 8'b00000110; 
    { 8'h6a, 4'h4 }: pattern = 8'b00000000; 
    { 8'h6a, 4'h5 }: pattern = 8'b00001110; 
    { 8'h6a, 4'h6 }: pattern = 8'b00000110; 
    { 8'h6a, 4'h7 }: pattern = 8'b00000110; 
    { 8'h6a, 4'h8 }: pattern = 8'b00000110; 
    { 8'h6a, 4'h9 }: pattern = 8'b00000110; 
    { 8'h6a, 4'ha }: pattern = 8'b00000110; 
    { 8'h6a, 4'hb }: pattern = 8'b00000110; 
    { 8'h6a, 4'hc }: pattern = 8'b01100110; 
    { 8'h6a, 4'hd }: pattern = 8'b01100110; 
    { 8'h6a, 4'he }: pattern = 8'b00111100; 
    { 8'h6a, 4'hf }: pattern = 8'b00000000; 

    { 8'h6b, 4'h0 }: pattern = 8'b00000000; 
    { 8'h6b, 4'h1 }: pattern = 8'b00000000; 
    { 8'h6b, 4'h2 }: pattern = 8'b11100000; 
    { 8'h6b, 4'h3 }: pattern = 8'b01100000; 
    { 8'h6b, 4'h4 }: pattern = 8'b01100000; 
    { 8'h6b, 4'h5 }: pattern = 8'b01100110; 
    { 8'h6b, 4'h6 }: pattern = 8'b01101100; 
    { 8'h6b, 4'h7 }: pattern = 8'b01111000; 
    { 8'h6b, 4'h8 }: pattern = 8'b01111000; 
    { 8'h6b, 4'h9 }: pattern = 8'b01101100; 
    { 8'h6b, 4'ha }: pattern = 8'b01100110; 
    { 8'h6b, 4'hb }: pattern = 8'b11100110; 
    { 8'h6b, 4'hc }: pattern = 8'b00000000; 
    { 8'h6b, 4'hd }: pattern = 8'b00000000; 
    { 8'h6b, 4'he }: pattern = 8'b00000000; 
    { 8'h6b, 4'hf }: pattern = 8'b00000000; 

    { 8'h6c, 4'h0 }: pattern = 8'b00000000; 
    { 8'h6c, 4'h1 }: pattern = 8'b00000000; 
    { 8'h6c, 4'h2 }: pattern = 8'b00111000; 
    { 8'h6c, 4'h3 }: pattern = 8'b00011000; 
    { 8'h6c, 4'h4 }: pattern = 8'b00011000; 
    { 8'h6c, 4'h5 }: pattern = 8'b00011000; 
    { 8'h6c, 4'h6 }: pattern = 8'b00011000; 
    { 8'h6c, 4'h7 }: pattern = 8'b00011000; 
    { 8'h6c, 4'h8 }: pattern = 8'b00011000; 
    { 8'h6c, 4'h9 }: pattern = 8'b00011000; 
    { 8'h6c, 4'ha }: pattern = 8'b00011000; 
    { 8'h6c, 4'hb }: pattern = 8'b00111100; 
    { 8'h6c, 4'hc }: pattern = 8'b00000000; 
    { 8'h6c, 4'hd }: pattern = 8'b00000000; 
    { 8'h6c, 4'he }: pattern = 8'b00000000; 
    { 8'h6c, 4'hf }: pattern = 8'b00000000; 

    { 8'h6d, 4'h0 }: pattern = 8'b00000000; 
    { 8'h6d, 4'h1 }: pattern = 8'b00000000; 
    { 8'h6d, 4'h2 }: pattern = 8'b00000000; 
    { 8'h6d, 4'h3 }: pattern = 8'b00000000; 
    { 8'h6d, 4'h4 }: pattern = 8'b00000000; 
    { 8'h6d, 4'h5 }: pattern = 8'b11101100; 
    { 8'h6d, 4'h6 }: pattern = 8'b11111110; 
    { 8'h6d, 4'h7 }: pattern = 8'b11010110; 
    { 8'h6d, 4'h8 }: pattern = 8'b11010110; 
    { 8'h6d, 4'h9 }: pattern = 8'b11010110; 
    { 8'h6d, 4'ha }: pattern = 8'b11010110; 
    { 8'h6d, 4'hb }: pattern = 8'b11000110; 
    { 8'h6d, 4'hc }: pattern = 8'b00000000; 
    { 8'h6d, 4'hd }: pattern = 8'b00000000; 
    { 8'h6d, 4'he }: pattern = 8'b00000000; 
    { 8'h6d, 4'hf }: pattern = 8'b00000000; 

    { 8'h6e, 4'h0 }: pattern = 8'b00000000; 
    { 8'h6e, 4'h1 }: pattern = 8'b00000000; 
    { 8'h6e, 4'h2 }: pattern = 8'b00000000; 
    { 8'h6e, 4'h3 }: pattern = 8'b00000000; 
    { 8'h6e, 4'h4 }: pattern = 8'b00000000; 
    { 8'h6e, 4'h5 }: pattern = 8'b11011100; 
    { 8'h6e, 4'h6 }: pattern = 8'b01100110; 
    { 8'h6e, 4'h7 }: pattern = 8'b01100110; 
    { 8'h6e, 4'h8 }: pattern = 8'b01100110; 
    { 8'h6e, 4'h9 }: pattern = 8'b01100110; 
    { 8'h6e, 4'ha }: pattern = 8'b01100110; 
    { 8'h6e, 4'hb }: pattern = 8'b01100110; 
    { 8'h6e, 4'hc }: pattern = 8'b00000000; 
    { 8'h6e, 4'hd }: pattern = 8'b00000000; 
    { 8'h6e, 4'he }: pattern = 8'b00000000; 
    { 8'h6e, 4'hf }: pattern = 8'b00000000; 

    { 8'h6f, 4'h0 }: pattern = 8'b00000000; 
    { 8'h6f, 4'h1 }: pattern = 8'b00000000; 
    { 8'h6f, 4'h2 }: pattern = 8'b00000000; 
    { 8'h6f, 4'h3 }: pattern = 8'b00000000; 
    { 8'h6f, 4'h4 }: pattern = 8'b00000000; 
    { 8'h6f, 4'h5 }: pattern = 8'b01111100; 
    { 8'h6f, 4'h6 }: pattern = 8'b11000110; 
    { 8'h6f, 4'h7 }: pattern = 8'b11000110; 
    { 8'h6f, 4'h8 }: pattern = 8'b11000110; 
    { 8'h6f, 4'h9 }: pattern = 8'b11000110; 
    { 8'h6f, 4'ha }: pattern = 8'b11000110; 
    { 8'h6f, 4'hb }: pattern = 8'b01111100; 
    { 8'h6f, 4'hc }: pattern = 8'b00000000; 
    { 8'h6f, 4'hd }: pattern = 8'b00000000; 
    { 8'h6f, 4'he }: pattern = 8'b00000000; 
    { 8'h6f, 4'hf }: pattern = 8'b00000000; 

    { 8'h70, 4'h0 }: pattern = 8'b00000000; 
    { 8'h70, 4'h1 }: pattern = 8'b00000000; 
    { 8'h70, 4'h2 }: pattern = 8'b00000000; 
    { 8'h70, 4'h3 }: pattern = 8'b00000000; 
    { 8'h70, 4'h4 }: pattern = 8'b00000000; 
    { 8'h70, 4'h5 }: pattern = 8'b11011100; 
    { 8'h70, 4'h6 }: pattern = 8'b01100110; 
    { 8'h70, 4'h7 }: pattern = 8'b01100110; 
    { 8'h70, 4'h8 }: pattern = 8'b01100110; 
    { 8'h70, 4'h9 }: pattern = 8'b01100110; 
    { 8'h70, 4'ha }: pattern = 8'b01100110; 
    { 8'h70, 4'hb }: pattern = 8'b01111100; 
    { 8'h70, 4'hc }: pattern = 8'b01100000; 
    { 8'h70, 4'hd }: pattern = 8'b01100000; 
    { 8'h70, 4'he }: pattern = 8'b11110000; 
    { 8'h70, 4'hf }: pattern = 8'b00000000; 

    { 8'h71, 4'h0 }: pattern = 8'b00000000; 
    { 8'h71, 4'h1 }: pattern = 8'b00000000; 
    { 8'h71, 4'h2 }: pattern = 8'b00000000; 
    { 8'h71, 4'h3 }: pattern = 8'b00000000; 
    { 8'h71, 4'h4 }: pattern = 8'b00000000; 
    { 8'h71, 4'h5 }: pattern = 8'b01110110; 
    { 8'h71, 4'h6 }: pattern = 8'b11001100; 
    { 8'h71, 4'h7 }: pattern = 8'b11001100; 
    { 8'h71, 4'h8 }: pattern = 8'b11001100; 
    { 8'h71, 4'h9 }: pattern = 8'b11001100; 
    { 8'h71, 4'ha }: pattern = 8'b11001100; 
    { 8'h71, 4'hb }: pattern = 8'b01111100; 
    { 8'h71, 4'hc }: pattern = 8'b00001100; 
    { 8'h71, 4'hd }: pattern = 8'b00001100; 
    { 8'h71, 4'he }: pattern = 8'b00011110; 
    { 8'h71, 4'hf }: pattern = 8'b00000000; 

    { 8'h72, 4'h0 }: pattern = 8'b00000000; 
    { 8'h72, 4'h1 }: pattern = 8'b00000000; 
    { 8'h72, 4'h2 }: pattern = 8'b00000000; 
    { 8'h72, 4'h3 }: pattern = 8'b00000000; 
    { 8'h72, 4'h4 }: pattern = 8'b00000000; 
    { 8'h72, 4'h5 }: pattern = 8'b11011100; 
    { 8'h72, 4'h6 }: pattern = 8'b01110110; 
    { 8'h72, 4'h7 }: pattern = 8'b01100110; 
    { 8'h72, 4'h8 }: pattern = 8'b01100000; 
    { 8'h72, 4'h9 }: pattern = 8'b01100000; 
    { 8'h72, 4'ha }: pattern = 8'b01100000; 
    { 8'h72, 4'hb }: pattern = 8'b11110000; 
    { 8'h72, 4'hc }: pattern = 8'b00000000; 
    { 8'h72, 4'hd }: pattern = 8'b00000000; 
    { 8'h72, 4'he }: pattern = 8'b00000000; 
    { 8'h72, 4'hf }: pattern = 8'b00000000; 

    { 8'h73, 4'h0 }: pattern = 8'b00000000; 
    { 8'h73, 4'h1 }: pattern = 8'b00000000; 
    { 8'h73, 4'h2 }: pattern = 8'b00000000; 
    { 8'h73, 4'h3 }: pattern = 8'b00000000; 
    { 8'h73, 4'h4 }: pattern = 8'b00000000; 
    { 8'h73, 4'h5 }: pattern = 8'b01111100; 
    { 8'h73, 4'h6 }: pattern = 8'b11000110; 
    { 8'h73, 4'h7 }: pattern = 8'b01100000; 
    { 8'h73, 4'h8 }: pattern = 8'b00111000; 
    { 8'h73, 4'h9 }: pattern = 8'b00001100; 
    { 8'h73, 4'ha }: pattern = 8'b11000110; 
    { 8'h73, 4'hb }: pattern = 8'b01111100; 
    { 8'h73, 4'hc }: pattern = 8'b00000000; 
    { 8'h73, 4'hd }: pattern = 8'b00000000; 
    { 8'h73, 4'he }: pattern = 8'b00000000; 
    { 8'h73, 4'hf }: pattern = 8'b00000000; 

    { 8'h74, 4'h0 }: pattern = 8'b00000000; 
    { 8'h74, 4'h1 }: pattern = 8'b00000000; 
    { 8'h74, 4'h2 }: pattern = 8'b00010000; 
    { 8'h74, 4'h3 }: pattern = 8'b00110000; 
    { 8'h74, 4'h4 }: pattern = 8'b00110000; 
    { 8'h74, 4'h5 }: pattern = 8'b11111100; 
    { 8'h74, 4'h6 }: pattern = 8'b00110000; 
    { 8'h74, 4'h7 }: pattern = 8'b00110000; 
    { 8'h74, 4'h8 }: pattern = 8'b00110000; 
    { 8'h74, 4'h9 }: pattern = 8'b00110000; 
    { 8'h74, 4'ha }: pattern = 8'b00110110; 
    { 8'h74, 4'hb }: pattern = 8'b00011100; 
    { 8'h74, 4'hc }: pattern = 8'b00000000; 
    { 8'h74, 4'hd }: pattern = 8'b00000000; 
    { 8'h74, 4'he }: pattern = 8'b00000000; 
    { 8'h74, 4'hf }: pattern = 8'b00000000; 

    { 8'h75, 4'h0 }: pattern = 8'b00000000; 
    { 8'h75, 4'h1 }: pattern = 8'b00000000; 
    { 8'h75, 4'h2 }: pattern = 8'b00000000; 
    { 8'h75, 4'h3 }: pattern = 8'b00000000; 
    { 8'h75, 4'h4 }: pattern = 8'b00000000; 
    { 8'h75, 4'h5 }: pattern = 8'b11001100; 
    { 8'h75, 4'h6 }: pattern = 8'b11001100; 
    { 8'h75, 4'h7 }: pattern = 8'b11001100; 
    { 8'h75, 4'h8 }: pattern = 8'b11001100; 
    { 8'h75, 4'h9 }: pattern = 8'b11001100; 
    { 8'h75, 4'ha }: pattern = 8'b11001100; 
    { 8'h75, 4'hb }: pattern = 8'b01110110; 
    { 8'h75, 4'hc }: pattern = 8'b00000000; 
    { 8'h75, 4'hd }: pattern = 8'b00000000; 
    { 8'h75, 4'he }: pattern = 8'b00000000; 
    { 8'h75, 4'hf }: pattern = 8'b00000000; 

    { 8'h76, 4'h0 }: pattern = 8'b00000000; 
    { 8'h76, 4'h1 }: pattern = 8'b00000000; 
    { 8'h76, 4'h2 }: pattern = 8'b00000000; 
    { 8'h76, 4'h3 }: pattern = 8'b00000000; 
    { 8'h76, 4'h4 }: pattern = 8'b00000000; 
    { 8'h76, 4'h5 }: pattern = 8'b01100110; 
    { 8'h76, 4'h6 }: pattern = 8'b01100110; 
    { 8'h76, 4'h7 }: pattern = 8'b01100110; 
    { 8'h76, 4'h8 }: pattern = 8'b01100110; 
    { 8'h76, 4'h9 }: pattern = 8'b01100110; 
    { 8'h76, 4'ha }: pattern = 8'b00111100; 
    { 8'h76, 4'hb }: pattern = 8'b00011000; 
    { 8'h76, 4'hc }: pattern = 8'b00000000; 
    { 8'h76, 4'hd }: pattern = 8'b00000000; 
    { 8'h76, 4'he }: pattern = 8'b00000000; 
    { 8'h76, 4'hf }: pattern = 8'b00000000; 

    { 8'h77, 4'h0 }: pattern = 8'b00000000; 
    { 8'h77, 4'h1 }: pattern = 8'b00000000; 
    { 8'h77, 4'h2 }: pattern = 8'b00000000; 
    { 8'h77, 4'h3 }: pattern = 8'b00000000; 
    { 8'h77, 4'h4 }: pattern = 8'b00000000; 
    { 8'h77, 4'h5 }: pattern = 8'b11000110; 
    { 8'h77, 4'h6 }: pattern = 8'b11000110; 
    { 8'h77, 4'h7 }: pattern = 8'b11010110; 
    { 8'h77, 4'h8 }: pattern = 8'b11010110; 
    { 8'h77, 4'h9 }: pattern = 8'b11010110; 
    { 8'h77, 4'ha }: pattern = 8'b11111110; 
    { 8'h77, 4'hb }: pattern = 8'b01101100; 
    { 8'h77, 4'hc }: pattern = 8'b00000000; 
    { 8'h77, 4'hd }: pattern = 8'b00000000; 
    { 8'h77, 4'he }: pattern = 8'b00000000; 
    { 8'h77, 4'hf }: pattern = 8'b00000000; 

    { 8'h78, 4'h0 }: pattern = 8'b00000000; 
    { 8'h78, 4'h1 }: pattern = 8'b00000000; 
    { 8'h78, 4'h2 }: pattern = 8'b00000000; 
    { 8'h78, 4'h3 }: pattern = 8'b00000000; 
    { 8'h78, 4'h4 }: pattern = 8'b00000000; 
    { 8'h78, 4'h5 }: pattern = 8'b11000110; 
    { 8'h78, 4'h6 }: pattern = 8'b01101100; 
    { 8'h78, 4'h7 }: pattern = 8'b00111000; 
    { 8'h78, 4'h8 }: pattern = 8'b00111000; 
    { 8'h78, 4'h9 }: pattern = 8'b00111000; 
    { 8'h78, 4'ha }: pattern = 8'b01101100; 
    { 8'h78, 4'hb }: pattern = 8'b11000110; 
    { 8'h78, 4'hc }: pattern = 8'b00000000; 
    { 8'h78, 4'hd }: pattern = 8'b00000000; 
    { 8'h78, 4'he }: pattern = 8'b00000000; 
    { 8'h78, 4'hf }: pattern = 8'b00000000; 

    { 8'h79, 4'h0 }: pattern = 8'b00000000; 
    { 8'h79, 4'h1 }: pattern = 8'b00000000; 
    { 8'h79, 4'h2 }: pattern = 8'b00000000; 
    { 8'h79, 4'h3 }: pattern = 8'b00000000; 
    { 8'h79, 4'h4 }: pattern = 8'b00000000; 
    { 8'h79, 4'h5 }: pattern = 8'b11000110; 
    { 8'h79, 4'h6 }: pattern = 8'b11000110; 
    { 8'h79, 4'h7 }: pattern = 8'b11000110; 
    { 8'h79, 4'h8 }: pattern = 8'b11000110; 
    { 8'h79, 4'h9 }: pattern = 8'b11000110; 
    { 8'h79, 4'ha }: pattern = 8'b11000110; 
    { 8'h79, 4'hb }: pattern = 8'b01111110; 
    { 8'h79, 4'hc }: pattern = 8'b00000110; 
    { 8'h79, 4'hd }: pattern = 8'b00001100; 
    { 8'h79, 4'he }: pattern = 8'b11111000; 
    { 8'h79, 4'hf }: pattern = 8'b00000000; 

    { 8'h7a, 4'h0 }: pattern = 8'b00000000; 
    { 8'h7a, 4'h1 }: pattern = 8'b00000000; 
    { 8'h7a, 4'h2 }: pattern = 8'b00000000; 
    { 8'h7a, 4'h3 }: pattern = 8'b00000000; 
    { 8'h7a, 4'h4 }: pattern = 8'b00000000; 
    { 8'h7a, 4'h5 }: pattern = 8'b11111110; 
    { 8'h7a, 4'h6 }: pattern = 8'b11001100; 
    { 8'h7a, 4'h7 }: pattern = 8'b00011000; 
    { 8'h7a, 4'h8 }: pattern = 8'b00110000; 
    { 8'h7a, 4'h9 }: pattern = 8'b01100000; 
    { 8'h7a, 4'ha }: pattern = 8'b11000110; 
    { 8'h7a, 4'hb }: pattern = 8'b11111110; 
    { 8'h7a, 4'hc }: pattern = 8'b00000000; 
    { 8'h7a, 4'hd }: pattern = 8'b00000000; 
    { 8'h7a, 4'he }: pattern = 8'b00000000; 
    { 8'h7a, 4'hf }: pattern = 8'b00000000; 

    { 8'h7b, 4'h0 }: pattern = 8'b00000000; 
    { 8'h7b, 4'h1 }: pattern = 8'b00000000; 
    { 8'h7b, 4'h2 }: pattern = 8'b00001110; 
    { 8'h7b, 4'h3 }: pattern = 8'b00011000; 
    { 8'h7b, 4'h4 }: pattern = 8'b00011000; 
    { 8'h7b, 4'h5 }: pattern = 8'b00011000; 
    { 8'h7b, 4'h6 }: pattern = 8'b01110000; 
    { 8'h7b, 4'h7 }: pattern = 8'b00011000; 
    { 8'h7b, 4'h8 }: pattern = 8'b00011000; 
    { 8'h7b, 4'h9 }: pattern = 8'b00011000; 
    { 8'h7b, 4'ha }: pattern = 8'b00011000; 
    { 8'h7b, 4'hb }: pattern = 8'b00001110; 
    { 8'h7b, 4'hc }: pattern = 8'b00000000; 
    { 8'h7b, 4'hd }: pattern = 8'b00000000; 
    { 8'h7b, 4'he }: pattern = 8'b00000000; 
    { 8'h7b, 4'hf }: pattern = 8'b00000000; 

    { 8'h7c, 4'h0 }: pattern = 8'b00000000; 
    { 8'h7c, 4'h1 }: pattern = 8'b00000000; 
    { 8'h7c, 4'h2 }: pattern = 8'b00011000; 
    { 8'h7c, 4'h3 }: pattern = 8'b00011000; 
    { 8'h7c, 4'h4 }: pattern = 8'b00011000; 
    { 8'h7c, 4'h5 }: pattern = 8'b00011000; 
    { 8'h7c, 4'h6 }: pattern = 8'b00000000; 
    { 8'h7c, 4'h7 }: pattern = 8'b00011000; 
    { 8'h7c, 4'h8 }: pattern = 8'b00011000; 
    { 8'h7c, 4'h9 }: pattern = 8'b00011000; 
    { 8'h7c, 4'ha }: pattern = 8'b00011000; 
    { 8'h7c, 4'hb }: pattern = 8'b00011000; 
    { 8'h7c, 4'hc }: pattern = 8'b00000000; 
    { 8'h7c, 4'hd }: pattern = 8'b00000000; 
    { 8'h7c, 4'he }: pattern = 8'b00000000; 
    { 8'h7c, 4'hf }: pattern = 8'b00000000; 

    { 8'h7d, 4'h0 }: pattern = 8'b00000000; 
    { 8'h7d, 4'h1 }: pattern = 8'b00000000; 
    { 8'h7d, 4'h2 }: pattern = 8'b01110000; 
    { 8'h7d, 4'h3 }: pattern = 8'b00011000; 
    { 8'h7d, 4'h4 }: pattern = 8'b00011000; 
    { 8'h7d, 4'h5 }: pattern = 8'b00011000; 
    { 8'h7d, 4'h6 }: pattern = 8'b00001110; 
    { 8'h7d, 4'h7 }: pattern = 8'b00011000; 
    { 8'h7d, 4'h8 }: pattern = 8'b00011000; 
    { 8'h7d, 4'h9 }: pattern = 8'b00011000; 
    { 8'h7d, 4'ha }: pattern = 8'b00011000; 
    { 8'h7d, 4'hb }: pattern = 8'b01110000; 
    { 8'h7d, 4'hc }: pattern = 8'b00000000; 
    { 8'h7d, 4'hd }: pattern = 8'b00000000; 
    { 8'h7d, 4'he }: pattern = 8'b00000000; 
    { 8'h7d, 4'hf }: pattern = 8'b00000000; 

    { 8'h7e, 4'h0 }: pattern = 8'b00000000; 
    { 8'h7e, 4'h1 }: pattern = 8'b00000000; 
    { 8'h7e, 4'h2 }: pattern = 8'b01110110; 
    { 8'h7e, 4'h3 }: pattern = 8'b11011100; 
    { 8'h7e, 4'h4 }: pattern = 8'b00000000; 
    { 8'h7e, 4'h5 }: pattern = 8'b00000000; 
    { 8'h7e, 4'h6 }: pattern = 8'b00000000; 
    { 8'h7e, 4'h7 }: pattern = 8'b00000000; 
    { 8'h7e, 4'h8 }: pattern = 8'b00000000; 
    { 8'h7e, 4'h9 }: pattern = 8'b00000000; 
    { 8'h7e, 4'ha }: pattern = 8'b00000000; 
    { 8'h7e, 4'hb }: pattern = 8'b00000000; 
    { 8'h7e, 4'hc }: pattern = 8'b00000000; 
    { 8'h7e, 4'hd }: pattern = 8'b00000000; 
    { 8'h7e, 4'he }: pattern = 8'b00000000; 
    { 8'h7e, 4'hf }: pattern = 8'b00000000; 

    { 8'h7f, 4'h0 }: pattern = 8'b00000000; 
    { 8'h7f, 4'h1 }: pattern = 8'b00000000; 
    { 8'h7f, 4'h2 }: pattern = 8'b00000000; 
    { 8'h7f, 4'h3 }: pattern = 8'b00000000; 
    { 8'h7f, 4'h4 }: pattern = 8'b00010000; 
    { 8'h7f, 4'h5 }: pattern = 8'b00111000; 
    { 8'h7f, 4'h6 }: pattern = 8'b01101100; 
    { 8'h7f, 4'h7 }: pattern = 8'b11000110; 
    { 8'h7f, 4'h8 }: pattern = 8'b11000110; 
    { 8'h7f, 4'h9 }: pattern = 8'b11000110; 
    { 8'h7f, 4'ha }: pattern = 8'b11111110; 
    { 8'h7f, 4'hb }: pattern = 8'b00000000; 
    { 8'h7f, 4'hc }: pattern = 8'b00000000; 
    { 8'h7f, 4'hd }: pattern = 8'b00000000; 
    { 8'h7f, 4'he }: pattern = 8'b00000000; 
    { 8'h7f, 4'hf }: pattern = 8'b00000000; 

    { 8'h80, 4'h0 }: pattern = 8'b00000000; 
    { 8'h80, 4'h1 }: pattern = 8'b00000000; 
    { 8'h80, 4'h2 }: pattern = 8'b00111100; 
    { 8'h80, 4'h3 }: pattern = 8'b01100110; 
    { 8'h80, 4'h4 }: pattern = 8'b11000010; 
    { 8'h80, 4'h5 }: pattern = 8'b11000000; 
    { 8'h80, 4'h6 }: pattern = 8'b11000000; 
    { 8'h80, 4'h7 }: pattern = 8'b11000000; 
    { 8'h80, 4'h8 }: pattern = 8'b11000010; 
    { 8'h80, 4'h9 }: pattern = 8'b01100110; 
    { 8'h80, 4'ha }: pattern = 8'b00111100; 
    { 8'h80, 4'hb }: pattern = 8'b00001100; 
    { 8'h80, 4'hc }: pattern = 8'b00000110; 
    { 8'h80, 4'hd }: pattern = 8'b01111100; 
    { 8'h80, 4'he }: pattern = 8'b00000000; 
    { 8'h80, 4'hf }: pattern = 8'b00000000; 

    { 8'h81, 4'h0 }: pattern = 8'b00000000; 
    { 8'h81, 4'h1 }: pattern = 8'b00000000; 
    { 8'h81, 4'h2 }: pattern = 8'b11001100; 
    { 8'h81, 4'h3 }: pattern = 8'b00000000; 
    { 8'h81, 4'h4 }: pattern = 8'b00000000; 
    { 8'h81, 4'h5 }: pattern = 8'b11001100; 
    { 8'h81, 4'h6 }: pattern = 8'b11001100; 
    { 8'h81, 4'h7 }: pattern = 8'b11001100; 
    { 8'h81, 4'h8 }: pattern = 8'b11001100; 
    { 8'h81, 4'h9 }: pattern = 8'b11001100; 
    { 8'h81, 4'ha }: pattern = 8'b11001100; 
    { 8'h81, 4'hb }: pattern = 8'b01110110; 
    { 8'h81, 4'hc }: pattern = 8'b00000000; 
    { 8'h81, 4'hd }: pattern = 8'b00000000; 
    { 8'h81, 4'he }: pattern = 8'b00000000; 
    { 8'h81, 4'hf }: pattern = 8'b00000000; 

    { 8'h82, 4'h0 }: pattern = 8'b00000000; 
    { 8'h82, 4'h1 }: pattern = 8'b00001100; 
    { 8'h82, 4'h2 }: pattern = 8'b00011000; 
    { 8'h82, 4'h3 }: pattern = 8'b00110000; 
    { 8'h82, 4'h4 }: pattern = 8'b00000000; 
    { 8'h82, 4'h5 }: pattern = 8'b01111100; 
    { 8'h82, 4'h6 }: pattern = 8'b11000110; 
    { 8'h82, 4'h7 }: pattern = 8'b11111110; 
    { 8'h82, 4'h8 }: pattern = 8'b11000000; 
    { 8'h82, 4'h9 }: pattern = 8'b11000000; 
    { 8'h82, 4'ha }: pattern = 8'b11000110; 
    { 8'h82, 4'hb }: pattern = 8'b01111100; 
    { 8'h82, 4'hc }: pattern = 8'b00000000; 
    { 8'h82, 4'hd }: pattern = 8'b00000000; 
    { 8'h82, 4'he }: pattern = 8'b00000000; 
    { 8'h82, 4'hf }: pattern = 8'b00000000; 

    { 8'h83, 4'h0 }: pattern = 8'b00000000; 
    { 8'h83, 4'h1 }: pattern = 8'b00010000; 
    { 8'h83, 4'h2 }: pattern = 8'b00111000; 
    { 8'h83, 4'h3 }: pattern = 8'b01101100; 
    { 8'h83, 4'h4 }: pattern = 8'b00000000; 
    { 8'h83, 4'h5 }: pattern = 8'b01111000; 
    { 8'h83, 4'h6 }: pattern = 8'b00001100; 
    { 8'h83, 4'h7 }: pattern = 8'b01111100; 
    { 8'h83, 4'h8 }: pattern = 8'b11001100; 
    { 8'h83, 4'h9 }: pattern = 8'b11001100; 
    { 8'h83, 4'ha }: pattern = 8'b11001100; 
    { 8'h83, 4'hb }: pattern = 8'b01110110; 
    { 8'h83, 4'hc }: pattern = 8'b00000000; 
    { 8'h83, 4'hd }: pattern = 8'b00000000; 
    { 8'h83, 4'he }: pattern = 8'b00000000; 
    { 8'h83, 4'hf }: pattern = 8'b00000000; 

    { 8'h84, 4'h0 }: pattern = 8'b00000000; 
    { 8'h84, 4'h1 }: pattern = 8'b00000000; 
    { 8'h84, 4'h2 }: pattern = 8'b11001100; 
    { 8'h84, 4'h3 }: pattern = 8'b00000000; 
    { 8'h84, 4'h4 }: pattern = 8'b00000000; 
    { 8'h84, 4'h5 }: pattern = 8'b01111000; 
    { 8'h84, 4'h6 }: pattern = 8'b00001100; 
    { 8'h84, 4'h7 }: pattern = 8'b01111100; 
    { 8'h84, 4'h8 }: pattern = 8'b11001100; 
    { 8'h84, 4'h9 }: pattern = 8'b11001100; 
    { 8'h84, 4'ha }: pattern = 8'b11001100; 
    { 8'h84, 4'hb }: pattern = 8'b01110110; 
    { 8'h84, 4'hc }: pattern = 8'b00000000; 
    { 8'h84, 4'hd }: pattern = 8'b00000000; 
    { 8'h84, 4'he }: pattern = 8'b00000000; 
    { 8'h84, 4'hf }: pattern = 8'b00000000; 

    { 8'h85, 4'h0 }: pattern = 8'b00000000; 
    { 8'h85, 4'h1 }: pattern = 8'b01100000; 
    { 8'h85, 4'h2 }: pattern = 8'b00110000; 
    { 8'h85, 4'h3 }: pattern = 8'b00011000; 
    { 8'h85, 4'h4 }: pattern = 8'b00000000; 
    { 8'h85, 4'h5 }: pattern = 8'b01111000; 
    { 8'h85, 4'h6 }: pattern = 8'b00001100; 
    { 8'h85, 4'h7 }: pattern = 8'b01111100; 
    { 8'h85, 4'h8 }: pattern = 8'b11001100; 
    { 8'h85, 4'h9 }: pattern = 8'b11001100; 
    { 8'h85, 4'ha }: pattern = 8'b11001100; 
    { 8'h85, 4'hb }: pattern = 8'b01110110; 
    { 8'h85, 4'hc }: pattern = 8'b00000000; 
    { 8'h85, 4'hd }: pattern = 8'b00000000; 
    { 8'h85, 4'he }: pattern = 8'b00000000; 
    { 8'h85, 4'hf }: pattern = 8'b00000000; 

    { 8'h86, 4'h0 }: pattern = 8'b00000000; 
    { 8'h86, 4'h1 }: pattern = 8'b00111000; 
    { 8'h86, 4'h2 }: pattern = 8'b01101100; 
    { 8'h86, 4'h3 }: pattern = 8'b00111000; 
    { 8'h86, 4'h4 }: pattern = 8'b00000000; 
    { 8'h86, 4'h5 }: pattern = 8'b01111000; 
    { 8'h86, 4'h6 }: pattern = 8'b00001100; 
    { 8'h86, 4'h7 }: pattern = 8'b01111100; 
    { 8'h86, 4'h8 }: pattern = 8'b11001100; 
    { 8'h86, 4'h9 }: pattern = 8'b11001100; 
    { 8'h86, 4'ha }: pattern = 8'b11001100; 
    { 8'h86, 4'hb }: pattern = 8'b01110110; 
    { 8'h86, 4'hc }: pattern = 8'b00000000; 
    { 8'h86, 4'hd }: pattern = 8'b00000000; 
    { 8'h86, 4'he }: pattern = 8'b00000000; 
    { 8'h86, 4'hf }: pattern = 8'b00000000; 

    { 8'h87, 4'h0 }: pattern = 8'b00000000; 
    { 8'h87, 4'h1 }: pattern = 8'b00000000; 
    { 8'h87, 4'h2 }: pattern = 8'b00000000; 
    { 8'h87, 4'h3 }: pattern = 8'b00000000; 
    { 8'h87, 4'h4 }: pattern = 8'b00111100; 
    { 8'h87, 4'h5 }: pattern = 8'b01100110; 
    { 8'h87, 4'h6 }: pattern = 8'b01100000; 
    { 8'h87, 4'h7 }: pattern = 8'b01100000; 
    { 8'h87, 4'h8 }: pattern = 8'b01100110; 
    { 8'h87, 4'h9 }: pattern = 8'b00111100; 
    { 8'h87, 4'ha }: pattern = 8'b00001100; 
    { 8'h87, 4'hb }: pattern = 8'b00000110; 
    { 8'h87, 4'hc }: pattern = 8'b00111100; 
    { 8'h87, 4'hd }: pattern = 8'b00000000; 
    { 8'h87, 4'he }: pattern = 8'b00000000; 
    { 8'h87, 4'hf }: pattern = 8'b00000000; 

    { 8'h88, 4'h0 }: pattern = 8'b00000000; 
    { 8'h88, 4'h1 }: pattern = 8'b00010000; 
    { 8'h88, 4'h2 }: pattern = 8'b00111000; 
    { 8'h88, 4'h3 }: pattern = 8'b01101100; 
    { 8'h88, 4'h4 }: pattern = 8'b00000000; 
    { 8'h88, 4'h5 }: pattern = 8'b01111100; 
    { 8'h88, 4'h6 }: pattern = 8'b11000110; 
    { 8'h88, 4'h7 }: pattern = 8'b11111110; 
    { 8'h88, 4'h8 }: pattern = 8'b11000000; 
    { 8'h88, 4'h9 }: pattern = 8'b11000000; 
    { 8'h88, 4'ha }: pattern = 8'b11000110; 
    { 8'h88, 4'hb }: pattern = 8'b01111100; 
    { 8'h88, 4'hc }: pattern = 8'b00000000; 
    { 8'h88, 4'hd }: pattern = 8'b00000000; 
    { 8'h88, 4'he }: pattern = 8'b00000000; 
    { 8'h88, 4'hf }: pattern = 8'b00000000; 

    { 8'h89, 4'h0 }: pattern = 8'b00000000; 
    { 8'h89, 4'h1 }: pattern = 8'b00000000; 
    { 8'h89, 4'h2 }: pattern = 8'b11000110; 
    { 8'h89, 4'h3 }: pattern = 8'b00000000; 
    { 8'h89, 4'h4 }: pattern = 8'b00000000; 
    { 8'h89, 4'h5 }: pattern = 8'b01111100; 
    { 8'h89, 4'h6 }: pattern = 8'b11000110; 
    { 8'h89, 4'h7 }: pattern = 8'b11111110; 
    { 8'h89, 4'h8 }: pattern = 8'b11000000; 
    { 8'h89, 4'h9 }: pattern = 8'b11000000; 
    { 8'h89, 4'ha }: pattern = 8'b11000110; 
    { 8'h89, 4'hb }: pattern = 8'b01111100; 
    { 8'h89, 4'hc }: pattern = 8'b00000000; 
    { 8'h89, 4'hd }: pattern = 8'b00000000; 
    { 8'h89, 4'he }: pattern = 8'b00000000; 
    { 8'h89, 4'hf }: pattern = 8'b00000000; 

    { 8'h8a, 4'h0 }: pattern = 8'b00000000; 
    { 8'h8a, 4'h1 }: pattern = 8'b01100000; 
    { 8'h8a, 4'h2 }: pattern = 8'b00110000; 
    { 8'h8a, 4'h3 }: pattern = 8'b00011000; 
    { 8'h8a, 4'h4 }: pattern = 8'b00000000; 
    { 8'h8a, 4'h5 }: pattern = 8'b01111100; 
    { 8'h8a, 4'h6 }: pattern = 8'b11000110; 
    { 8'h8a, 4'h7 }: pattern = 8'b11111110; 
    { 8'h8a, 4'h8 }: pattern = 8'b11000000; 
    { 8'h8a, 4'h9 }: pattern = 8'b11000000; 
    { 8'h8a, 4'ha }: pattern = 8'b11000110; 
    { 8'h8a, 4'hb }: pattern = 8'b01111100; 
    { 8'h8a, 4'hc }: pattern = 8'b00000000; 
    { 8'h8a, 4'hd }: pattern = 8'b00000000; 
    { 8'h8a, 4'he }: pattern = 8'b00000000; 
    { 8'h8a, 4'hf }: pattern = 8'b00000000; 

    { 8'h8b, 4'h0 }: pattern = 8'b00000000; 
    { 8'h8b, 4'h1 }: pattern = 8'b00000000; 
    { 8'h8b, 4'h2 }: pattern = 8'b01100110; 
    { 8'h8b, 4'h3 }: pattern = 8'b00000000; 
    { 8'h8b, 4'h4 }: pattern = 8'b00000000; 
    { 8'h8b, 4'h5 }: pattern = 8'b00111000; 
    { 8'h8b, 4'h6 }: pattern = 8'b00011000; 
    { 8'h8b, 4'h7 }: pattern = 8'b00011000; 
    { 8'h8b, 4'h8 }: pattern = 8'b00011000; 
    { 8'h8b, 4'h9 }: pattern = 8'b00011000; 
    { 8'h8b, 4'ha }: pattern = 8'b00011000; 
    { 8'h8b, 4'hb }: pattern = 8'b00111100; 
    { 8'h8b, 4'hc }: pattern = 8'b00000000; 
    { 8'h8b, 4'hd }: pattern = 8'b00000000; 
    { 8'h8b, 4'he }: pattern = 8'b00000000; 
    { 8'h8b, 4'hf }: pattern = 8'b00000000; 

    { 8'h8c, 4'h0 }: pattern = 8'b00000000; 
    { 8'h8c, 4'h1 }: pattern = 8'b00011000; 
    { 8'h8c, 4'h2 }: pattern = 8'b00111100; 
    { 8'h8c, 4'h3 }: pattern = 8'b01100110; 
    { 8'h8c, 4'h4 }: pattern = 8'b00000000; 
    { 8'h8c, 4'h5 }: pattern = 8'b00111000; 
    { 8'h8c, 4'h6 }: pattern = 8'b00011000; 
    { 8'h8c, 4'h7 }: pattern = 8'b00011000; 
    { 8'h8c, 4'h8 }: pattern = 8'b00011000; 
    { 8'h8c, 4'h9 }: pattern = 8'b00011000; 
    { 8'h8c, 4'ha }: pattern = 8'b00011000; 
    { 8'h8c, 4'hb }: pattern = 8'b00111100; 
    { 8'h8c, 4'hc }: pattern = 8'b00000000; 
    { 8'h8c, 4'hd }: pattern = 8'b00000000; 
    { 8'h8c, 4'he }: pattern = 8'b00000000; 
    { 8'h8c, 4'hf }: pattern = 8'b00000000; 

    { 8'h8d, 4'h0 }: pattern = 8'b00000000; 
    { 8'h8d, 4'h1 }: pattern = 8'b01100000; 
    { 8'h8d, 4'h2 }: pattern = 8'b00110000; 
    { 8'h8d, 4'h3 }: pattern = 8'b00011000; 
    { 8'h8d, 4'h4 }: pattern = 8'b00000000; 
    { 8'h8d, 4'h5 }: pattern = 8'b00111000; 
    { 8'h8d, 4'h6 }: pattern = 8'b00011000; 
    { 8'h8d, 4'h7 }: pattern = 8'b00011000; 
    { 8'h8d, 4'h8 }: pattern = 8'b00011000; 
    { 8'h8d, 4'h9 }: pattern = 8'b00011000; 
    { 8'h8d, 4'ha }: pattern = 8'b00011000; 
    { 8'h8d, 4'hb }: pattern = 8'b00111100; 
    { 8'h8d, 4'hc }: pattern = 8'b00000000; 
    { 8'h8d, 4'hd }: pattern = 8'b00000000; 
    { 8'h8d, 4'he }: pattern = 8'b00000000; 
    { 8'h8d, 4'hf }: pattern = 8'b00000000; 

    { 8'h8e, 4'h0 }: pattern = 8'b00000000; 
    { 8'h8e, 4'h1 }: pattern = 8'b11000110; 
    { 8'h8e, 4'h2 }: pattern = 8'b00000000; 
    { 8'h8e, 4'h3 }: pattern = 8'b00010000; 
    { 8'h8e, 4'h4 }: pattern = 8'b00111000; 
    { 8'h8e, 4'h5 }: pattern = 8'b01101100; 
    { 8'h8e, 4'h6 }: pattern = 8'b11000110; 
    { 8'h8e, 4'h7 }: pattern = 8'b11000110; 
    { 8'h8e, 4'h8 }: pattern = 8'b11111110; 
    { 8'h8e, 4'h9 }: pattern = 8'b11000110; 
    { 8'h8e, 4'ha }: pattern = 8'b11000110; 
    { 8'h8e, 4'hb }: pattern = 8'b11000110; 
    { 8'h8e, 4'hc }: pattern = 8'b00000000; 
    { 8'h8e, 4'hd }: pattern = 8'b00000000; 
    { 8'h8e, 4'he }: pattern = 8'b00000000; 
    { 8'h8e, 4'hf }: pattern = 8'b00000000; 

    { 8'h8f, 4'h0 }: pattern = 8'b00111000; 
    { 8'h8f, 4'h1 }: pattern = 8'b01101100; 
    { 8'h8f, 4'h2 }: pattern = 8'b00111000; 
    { 8'h8f, 4'h3 }: pattern = 8'b00000000; 
    { 8'h8f, 4'h4 }: pattern = 8'b00111000; 
    { 8'h8f, 4'h5 }: pattern = 8'b01101100; 
    { 8'h8f, 4'h6 }: pattern = 8'b11000110; 
    { 8'h8f, 4'h7 }: pattern = 8'b11000110; 
    { 8'h8f, 4'h8 }: pattern = 8'b11111110; 
    { 8'h8f, 4'h9 }: pattern = 8'b11000110; 
    { 8'h8f, 4'ha }: pattern = 8'b11000110; 
    { 8'h8f, 4'hb }: pattern = 8'b11000110; 
    { 8'h8f, 4'hc }: pattern = 8'b00000000; 
    { 8'h8f, 4'hd }: pattern = 8'b00000000; 
    { 8'h8f, 4'he }: pattern = 8'b00000000; 
    { 8'h8f, 4'hf }: pattern = 8'b00000000; 

    { 8'h90, 4'h0 }: pattern = 8'b00011000; 
    { 8'h90, 4'h1 }: pattern = 8'b00110000; 
    { 8'h90, 4'h2 }: pattern = 8'b01100000; 
    { 8'h90, 4'h3 }: pattern = 8'b00000000; 
    { 8'h90, 4'h4 }: pattern = 8'b11111110; 
    { 8'h90, 4'h5 }: pattern = 8'b01100110; 
    { 8'h90, 4'h6 }: pattern = 8'b01100000; 
    { 8'h90, 4'h7 }: pattern = 8'b01111100; 
    { 8'h90, 4'h8 }: pattern = 8'b01100000; 
    { 8'h90, 4'h9 }: pattern = 8'b01100000; 
    { 8'h90, 4'ha }: pattern = 8'b01100110; 
    { 8'h90, 4'hb }: pattern = 8'b11111110; 
    { 8'h90, 4'hc }: pattern = 8'b00000000; 
    { 8'h90, 4'hd }: pattern = 8'b00000000; 
    { 8'h90, 4'he }: pattern = 8'b00000000; 
    { 8'h90, 4'hf }: pattern = 8'b00000000; 

    { 8'h91, 4'h0 }: pattern = 8'b00000000; 
    { 8'h91, 4'h1 }: pattern = 8'b00000000; 
    { 8'h91, 4'h2 }: pattern = 8'b00000000; 
    { 8'h91, 4'h3 }: pattern = 8'b00000000; 
    { 8'h91, 4'h4 }: pattern = 8'b00000000; 
    { 8'h91, 4'h5 }: pattern = 8'b11001100; 
    { 8'h91, 4'h6 }: pattern = 8'b01110110; 
    { 8'h91, 4'h7 }: pattern = 8'b00110110; 
    { 8'h91, 4'h8 }: pattern = 8'b01111110; 
    { 8'h91, 4'h9 }: pattern = 8'b11011000; 
    { 8'h91, 4'ha }: pattern = 8'b11011000; 
    { 8'h91, 4'hb }: pattern = 8'b01101110; 
    { 8'h91, 4'hc }: pattern = 8'b00000000; 
    { 8'h91, 4'hd }: pattern = 8'b00000000; 
    { 8'h91, 4'he }: pattern = 8'b00000000; 
    { 8'h91, 4'hf }: pattern = 8'b00000000; 

    { 8'h92, 4'h0 }: pattern = 8'b00000000; 
    { 8'h92, 4'h1 }: pattern = 8'b00000000; 
    { 8'h92, 4'h2 }: pattern = 8'b00111110; 
    { 8'h92, 4'h3 }: pattern = 8'b01101100; 
    { 8'h92, 4'h4 }: pattern = 8'b11001100; 
    { 8'h92, 4'h5 }: pattern = 8'b11001100; 
    { 8'h92, 4'h6 }: pattern = 8'b11111110; 
    { 8'h92, 4'h7 }: pattern = 8'b11001100; 
    { 8'h92, 4'h8 }: pattern = 8'b11001100; 
    { 8'h92, 4'h9 }: pattern = 8'b11001100; 
    { 8'h92, 4'ha }: pattern = 8'b11001100; 
    { 8'h92, 4'hb }: pattern = 8'b11001110; 
    { 8'h92, 4'hc }: pattern = 8'b00000000; 
    { 8'h92, 4'hd }: pattern = 8'b00000000; 
    { 8'h92, 4'he }: pattern = 8'b00000000; 
    { 8'h92, 4'hf }: pattern = 8'b00000000; 

    { 8'h93, 4'h0 }: pattern = 8'b00000000; 
    { 8'h93, 4'h1 }: pattern = 8'b00010000; 
    { 8'h93, 4'h2 }: pattern = 8'b00111000; 
    { 8'h93, 4'h3 }: pattern = 8'b01101100; 
    { 8'h93, 4'h4 }: pattern = 8'b00000000; 
    { 8'h93, 4'h5 }: pattern = 8'b01111100; 
    { 8'h93, 4'h6 }: pattern = 8'b11000110; 
    { 8'h93, 4'h7 }: pattern = 8'b11000110; 
    { 8'h93, 4'h8 }: pattern = 8'b11000110; 
    { 8'h93, 4'h9 }: pattern = 8'b11000110; 
    { 8'h93, 4'ha }: pattern = 8'b11000110; 
    { 8'h93, 4'hb }: pattern = 8'b01111100; 
    { 8'h93, 4'hc }: pattern = 8'b00000000; 
    { 8'h93, 4'hd }: pattern = 8'b00000000; 
    { 8'h93, 4'he }: pattern = 8'b00000000; 
    { 8'h93, 4'hf }: pattern = 8'b00000000; 

    { 8'h94, 4'h0 }: pattern = 8'b00000000; 
    { 8'h94, 4'h1 }: pattern = 8'b00000000; 
    { 8'h94, 4'h2 }: pattern = 8'b11000110; 
    { 8'h94, 4'h3 }: pattern = 8'b00000000; 
    { 8'h94, 4'h4 }: pattern = 8'b00000000; 
    { 8'h94, 4'h5 }: pattern = 8'b01111100; 
    { 8'h94, 4'h6 }: pattern = 8'b11000110; 
    { 8'h94, 4'h7 }: pattern = 8'b11000110; 
    { 8'h94, 4'h8 }: pattern = 8'b11000110; 
    { 8'h94, 4'h9 }: pattern = 8'b11000110; 
    { 8'h94, 4'ha }: pattern = 8'b11000110; 
    { 8'h94, 4'hb }: pattern = 8'b01111100; 
    { 8'h94, 4'hc }: pattern = 8'b00000000; 
    { 8'h94, 4'hd }: pattern = 8'b00000000; 
    { 8'h94, 4'he }: pattern = 8'b00000000; 
    { 8'h94, 4'hf }: pattern = 8'b00000000; 

    { 8'h95, 4'h0 }: pattern = 8'b00000000; 
    { 8'h95, 4'h1 }: pattern = 8'b01100000; 
    { 8'h95, 4'h2 }: pattern = 8'b00110000; 
    { 8'h95, 4'h3 }: pattern = 8'b00011000; 
    { 8'h95, 4'h4 }: pattern = 8'b00000000; 
    { 8'h95, 4'h5 }: pattern = 8'b01111100; 
    { 8'h95, 4'h6 }: pattern = 8'b11000110; 
    { 8'h95, 4'h7 }: pattern = 8'b11000110; 
    { 8'h95, 4'h8 }: pattern = 8'b11000110; 
    { 8'h95, 4'h9 }: pattern = 8'b11000110; 
    { 8'h95, 4'ha }: pattern = 8'b11000110; 
    { 8'h95, 4'hb }: pattern = 8'b01111100; 
    { 8'h95, 4'hc }: pattern = 8'b00000000; 
    { 8'h95, 4'hd }: pattern = 8'b00000000; 
    { 8'h95, 4'he }: pattern = 8'b00000000; 
    { 8'h95, 4'hf }: pattern = 8'b00000000; 

    { 8'h96, 4'h0 }: pattern = 8'b00000000; 
    { 8'h96, 4'h1 }: pattern = 8'b00110000; 
    { 8'h96, 4'h2 }: pattern = 8'b01111000; 
    { 8'h96, 4'h3 }: pattern = 8'b11001100; 
    { 8'h96, 4'h4 }: pattern = 8'b00000000; 
    { 8'h96, 4'h5 }: pattern = 8'b11001100; 
    { 8'h96, 4'h6 }: pattern = 8'b11001100; 
    { 8'h96, 4'h7 }: pattern = 8'b11001100; 
    { 8'h96, 4'h8 }: pattern = 8'b11001100; 
    { 8'h96, 4'h9 }: pattern = 8'b11001100; 
    { 8'h96, 4'ha }: pattern = 8'b11001100; 
    { 8'h96, 4'hb }: pattern = 8'b01110110; 
    { 8'h96, 4'hc }: pattern = 8'b00000000; 
    { 8'h96, 4'hd }: pattern = 8'b00000000; 
    { 8'h96, 4'he }: pattern = 8'b00000000; 
    { 8'h96, 4'hf }: pattern = 8'b00000000; 

    { 8'h97, 4'h0 }: pattern = 8'b00000000; 
    { 8'h97, 4'h1 }: pattern = 8'b01100000; 
    { 8'h97, 4'h2 }: pattern = 8'b00110000; 
    { 8'h97, 4'h3 }: pattern = 8'b00011000; 
    { 8'h97, 4'h4 }: pattern = 8'b00000000; 
    { 8'h97, 4'h5 }: pattern = 8'b11001100; 
    { 8'h97, 4'h6 }: pattern = 8'b11001100; 
    { 8'h97, 4'h7 }: pattern = 8'b11001100; 
    { 8'h97, 4'h8 }: pattern = 8'b11001100; 
    { 8'h97, 4'h9 }: pattern = 8'b11001100; 
    { 8'h97, 4'ha }: pattern = 8'b11001100; 
    { 8'h97, 4'hb }: pattern = 8'b01110110; 
    { 8'h97, 4'hc }: pattern = 8'b00000000; 
    { 8'h97, 4'hd }: pattern = 8'b00000000; 
    { 8'h97, 4'he }: pattern = 8'b00000000; 
    { 8'h97, 4'hf }: pattern = 8'b00000000; 

    { 8'h98, 4'h0 }: pattern = 8'b00000000; 
    { 8'h98, 4'h1 }: pattern = 8'b00000000; 
    { 8'h98, 4'h2 }: pattern = 8'b11000110; 
    { 8'h98, 4'h3 }: pattern = 8'b00000000; 
    { 8'h98, 4'h4 }: pattern = 8'b00000000; 
    { 8'h98, 4'h5 }: pattern = 8'b11000110; 
    { 8'h98, 4'h6 }: pattern = 8'b11000110; 
    { 8'h98, 4'h7 }: pattern = 8'b11000110; 
    { 8'h98, 4'h8 }: pattern = 8'b11000110; 
    { 8'h98, 4'h9 }: pattern = 8'b11000110; 
    { 8'h98, 4'ha }: pattern = 8'b11000110; 
    { 8'h98, 4'hb }: pattern = 8'b01111110; 
    { 8'h98, 4'hc }: pattern = 8'b00000110; 
    { 8'h98, 4'hd }: pattern = 8'b00001100; 
    { 8'h98, 4'he }: pattern = 8'b01111000; 
    { 8'h98, 4'hf }: pattern = 8'b00000000; 

    { 8'h99, 4'h0 }: pattern = 8'b00000000; 
    { 8'h99, 4'h1 }: pattern = 8'b11000110; 
    { 8'h99, 4'h2 }: pattern = 8'b00000000; 
    { 8'h99, 4'h3 }: pattern = 8'b01111100; 
    { 8'h99, 4'h4 }: pattern = 8'b11000110; 
    { 8'h99, 4'h5 }: pattern = 8'b11000110; 
    { 8'h99, 4'h6 }: pattern = 8'b11000110; 
    { 8'h99, 4'h7 }: pattern = 8'b11000110; 
    { 8'h99, 4'h8 }: pattern = 8'b11000110; 
    { 8'h99, 4'h9 }: pattern = 8'b11000110; 
    { 8'h99, 4'ha }: pattern = 8'b11000110; 
    { 8'h99, 4'hb }: pattern = 8'b01111100; 
    { 8'h99, 4'hc }: pattern = 8'b00000000; 
    { 8'h99, 4'hd }: pattern = 8'b00000000; 
    { 8'h99, 4'he }: pattern = 8'b00000000; 
    { 8'h99, 4'hf }: pattern = 8'b00000000; 

    { 8'h9a, 4'h0 }: pattern = 8'b00000000; 
    { 8'h9a, 4'h1 }: pattern = 8'b11000110; 
    { 8'h9a, 4'h2 }: pattern = 8'b00000000; 
    { 8'h9a, 4'h3 }: pattern = 8'b11000110; 
    { 8'h9a, 4'h4 }: pattern = 8'b11000110; 
    { 8'h9a, 4'h5 }: pattern = 8'b11000110; 
    { 8'h9a, 4'h6 }: pattern = 8'b11000110; 
    { 8'h9a, 4'h7 }: pattern = 8'b11000110; 
    { 8'h9a, 4'h8 }: pattern = 8'b11000110; 
    { 8'h9a, 4'h9 }: pattern = 8'b11000110; 
    { 8'h9a, 4'ha }: pattern = 8'b11000110; 
    { 8'h9a, 4'hb }: pattern = 8'b01111100; 
    { 8'h9a, 4'hc }: pattern = 8'b00000000; 
    { 8'h9a, 4'hd }: pattern = 8'b00000000; 
    { 8'h9a, 4'he }: pattern = 8'b00000000; 
    { 8'h9a, 4'hf }: pattern = 8'b00000000; 

    { 8'h9b, 4'h0 }: pattern = 8'b00000000; 
    { 8'h9b, 4'h1 }: pattern = 8'b00011000; 
    { 8'h9b, 4'h2 }: pattern = 8'b00011000; 
    { 8'h9b, 4'h3 }: pattern = 8'b00111100; 
    { 8'h9b, 4'h4 }: pattern = 8'b01100110; 
    { 8'h9b, 4'h5 }: pattern = 8'b01100000; 
    { 8'h9b, 4'h6 }: pattern = 8'b01100000; 
    { 8'h9b, 4'h7 }: pattern = 8'b01100000; 
    { 8'h9b, 4'h8 }: pattern = 8'b01100110; 
    { 8'h9b, 4'h9 }: pattern = 8'b00111100; 
    { 8'h9b, 4'ha }: pattern = 8'b00011000; 
    { 8'h9b, 4'hb }: pattern = 8'b00011000; 
    { 8'h9b, 4'hc }: pattern = 8'b00000000; 
    { 8'h9b, 4'hd }: pattern = 8'b00000000; 
    { 8'h9b, 4'he }: pattern = 8'b00000000; 
    { 8'h9b, 4'hf }: pattern = 8'b00000000; 

    { 8'h9c, 4'h0 }: pattern = 8'b00000000; 
    { 8'h9c, 4'h1 }: pattern = 8'b00111000; 
    { 8'h9c, 4'h2 }: pattern = 8'b01101100; 
    { 8'h9c, 4'h3 }: pattern = 8'b01100100; 
    { 8'h9c, 4'h4 }: pattern = 8'b01100000; 
    { 8'h9c, 4'h5 }: pattern = 8'b11110000; 
    { 8'h9c, 4'h6 }: pattern = 8'b01100000; 
    { 8'h9c, 4'h7 }: pattern = 8'b01100000; 
    { 8'h9c, 4'h8 }: pattern = 8'b01100000; 
    { 8'h9c, 4'h9 }: pattern = 8'b01100000; 
    { 8'h9c, 4'ha }: pattern = 8'b11100110; 
    { 8'h9c, 4'hb }: pattern = 8'b11111100; 
    { 8'h9c, 4'hc }: pattern = 8'b00000000; 
    { 8'h9c, 4'hd }: pattern = 8'b00000000; 
    { 8'h9c, 4'he }: pattern = 8'b00000000; 
    { 8'h9c, 4'hf }: pattern = 8'b00000000; 

    { 8'h9d, 4'h0 }: pattern = 8'b00000000; 
    { 8'h9d, 4'h1 }: pattern = 8'b00000000; 
    { 8'h9d, 4'h2 }: pattern = 8'b01100110; 
    { 8'h9d, 4'h3 }: pattern = 8'b01100110; 
    { 8'h9d, 4'h4 }: pattern = 8'b00111100; 
    { 8'h9d, 4'h5 }: pattern = 8'b00011000; 
    { 8'h9d, 4'h6 }: pattern = 8'b01111110; 
    { 8'h9d, 4'h7 }: pattern = 8'b00011000; 
    { 8'h9d, 4'h8 }: pattern = 8'b01111110; 
    { 8'h9d, 4'h9 }: pattern = 8'b00011000; 
    { 8'h9d, 4'ha }: pattern = 8'b00011000; 
    { 8'h9d, 4'hb }: pattern = 8'b00011000; 
    { 8'h9d, 4'hc }: pattern = 8'b00000000; 
    { 8'h9d, 4'hd }: pattern = 8'b00000000; 
    { 8'h9d, 4'he }: pattern = 8'b00000000; 
    { 8'h9d, 4'hf }: pattern = 8'b00000000; 

    { 8'h9e, 4'h0 }: pattern = 8'b00000000; 
    { 8'h9e, 4'h1 }: pattern = 8'b11111000; 
    { 8'h9e, 4'h2 }: pattern = 8'b11001100; 
    { 8'h9e, 4'h3 }: pattern = 8'b11001100; 
    { 8'h9e, 4'h4 }: pattern = 8'b11111000; 
    { 8'h9e, 4'h5 }: pattern = 8'b11000100; 
    { 8'h9e, 4'h6 }: pattern = 8'b11001100; 
    { 8'h9e, 4'h7 }: pattern = 8'b11011110; 
    { 8'h9e, 4'h8 }: pattern = 8'b11001100; 
    { 8'h9e, 4'h9 }: pattern = 8'b11001100; 
    { 8'h9e, 4'ha }: pattern = 8'b11001100; 
    { 8'h9e, 4'hb }: pattern = 8'b11000110; 
    { 8'h9e, 4'hc }: pattern = 8'b00000000; 
    { 8'h9e, 4'hd }: pattern = 8'b00000000; 
    { 8'h9e, 4'he }: pattern = 8'b00000000; 
    { 8'h9e, 4'hf }: pattern = 8'b00000000; 

    { 8'h9f, 4'h0 }: pattern = 8'b00000000; 
    { 8'h9f, 4'h1 }: pattern = 8'b00001110; 
    { 8'h9f, 4'h2 }: pattern = 8'b00011011; 
    { 8'h9f, 4'h3 }: pattern = 8'b00011000; 
    { 8'h9f, 4'h4 }: pattern = 8'b00011000; 
    { 8'h9f, 4'h5 }: pattern = 8'b00011000; 
    { 8'h9f, 4'h6 }: pattern = 8'b01111110; 
    { 8'h9f, 4'h7 }: pattern = 8'b00011000; 
    { 8'h9f, 4'h8 }: pattern = 8'b00011000; 
    { 8'h9f, 4'h9 }: pattern = 8'b00011000; 
    { 8'h9f, 4'ha }: pattern = 8'b00011000; 
    { 8'h9f, 4'hb }: pattern = 8'b00011000; 
    { 8'h9f, 4'hc }: pattern = 8'b11011000; 
    { 8'h9f, 4'hd }: pattern = 8'b01110000; 
    { 8'h9f, 4'he }: pattern = 8'b00000000; 
    { 8'h9f, 4'hf }: pattern = 8'b00000000; 

    { 8'ha0, 4'h0 }: pattern = 8'b00000000; 
    { 8'ha0, 4'h1 }: pattern = 8'b00011000; 
    { 8'ha0, 4'h2 }: pattern = 8'b00110000; 
    { 8'ha0, 4'h3 }: pattern = 8'b01100000; 
    { 8'ha0, 4'h4 }: pattern = 8'b00000000; 
    { 8'ha0, 4'h5 }: pattern = 8'b01111000; 
    { 8'ha0, 4'h6 }: pattern = 8'b00001100; 
    { 8'ha0, 4'h7 }: pattern = 8'b01111100; 
    { 8'ha0, 4'h8 }: pattern = 8'b11001100; 
    { 8'ha0, 4'h9 }: pattern = 8'b11001100; 
    { 8'ha0, 4'ha }: pattern = 8'b11001100; 
    { 8'ha0, 4'hb }: pattern = 8'b01110110; 
    { 8'ha0, 4'hc }: pattern = 8'b00000000; 
    { 8'ha0, 4'hd }: pattern = 8'b00000000; 
    { 8'ha0, 4'he }: pattern = 8'b00000000; 
    { 8'ha0, 4'hf }: pattern = 8'b00000000; 

    { 8'ha1, 4'h0 }: pattern = 8'b00000000; 
    { 8'ha1, 4'h1 }: pattern = 8'b00001100; 
    { 8'ha1, 4'h2 }: pattern = 8'b00011000; 
    { 8'ha1, 4'h3 }: pattern = 8'b00110000; 
    { 8'ha1, 4'h4 }: pattern = 8'b00000000; 
    { 8'ha1, 4'h5 }: pattern = 8'b00111000; 
    { 8'ha1, 4'h6 }: pattern = 8'b00011000; 
    { 8'ha1, 4'h7 }: pattern = 8'b00011000; 
    { 8'ha1, 4'h8 }: pattern = 8'b00011000; 
    { 8'ha1, 4'h9 }: pattern = 8'b00011000; 
    { 8'ha1, 4'ha }: pattern = 8'b00011000; 
    { 8'ha1, 4'hb }: pattern = 8'b00111100; 
    { 8'ha1, 4'hc }: pattern = 8'b00000000; 
    { 8'ha1, 4'hd }: pattern = 8'b00000000; 
    { 8'ha1, 4'he }: pattern = 8'b00000000; 
    { 8'ha1, 4'hf }: pattern = 8'b00000000; 

    { 8'ha2, 4'h0 }: pattern = 8'b00000000; 
    { 8'ha2, 4'h1 }: pattern = 8'b00011000; 
    { 8'ha2, 4'h2 }: pattern = 8'b00110000; 
    { 8'ha2, 4'h3 }: pattern = 8'b01100000; 
    { 8'ha2, 4'h4 }: pattern = 8'b00000000; 
    { 8'ha2, 4'h5 }: pattern = 8'b01111100; 
    { 8'ha2, 4'h6 }: pattern = 8'b11000110; 
    { 8'ha2, 4'h7 }: pattern = 8'b11000110; 
    { 8'ha2, 4'h8 }: pattern = 8'b11000110; 
    { 8'ha2, 4'h9 }: pattern = 8'b11000110; 
    { 8'ha2, 4'ha }: pattern = 8'b11000110; 
    { 8'ha2, 4'hb }: pattern = 8'b01111100; 
    { 8'ha2, 4'hc }: pattern = 8'b00000000; 
    { 8'ha2, 4'hd }: pattern = 8'b00000000; 
    { 8'ha2, 4'he }: pattern = 8'b00000000; 
    { 8'ha2, 4'hf }: pattern = 8'b00000000; 

    { 8'ha3, 4'h0 }: pattern = 8'b00000000; 
    { 8'ha3, 4'h1 }: pattern = 8'b00011000; 
    { 8'ha3, 4'h2 }: pattern = 8'b00110000; 
    { 8'ha3, 4'h3 }: pattern = 8'b01100000; 
    { 8'ha3, 4'h4 }: pattern = 8'b00000000; 
    { 8'ha3, 4'h5 }: pattern = 8'b11001100; 
    { 8'ha3, 4'h6 }: pattern = 8'b11001100; 
    { 8'ha3, 4'h7 }: pattern = 8'b11001100; 
    { 8'ha3, 4'h8 }: pattern = 8'b11001100; 
    { 8'ha3, 4'h9 }: pattern = 8'b11001100; 
    { 8'ha3, 4'ha }: pattern = 8'b11001100; 
    { 8'ha3, 4'hb }: pattern = 8'b01110110; 
    { 8'ha3, 4'hc }: pattern = 8'b00000000; 
    { 8'ha3, 4'hd }: pattern = 8'b00000000; 
    { 8'ha3, 4'he }: pattern = 8'b00000000; 
    { 8'ha3, 4'hf }: pattern = 8'b00000000; 

    { 8'ha4, 4'h0 }: pattern = 8'b00000000; 
    { 8'ha4, 4'h1 }: pattern = 8'b00000000; 
    { 8'ha4, 4'h2 }: pattern = 8'b01110110; 
    { 8'ha4, 4'h3 }: pattern = 8'b11011100; 
    { 8'ha4, 4'h4 }: pattern = 8'b00000000; 
    { 8'ha4, 4'h5 }: pattern = 8'b11011100; 
    { 8'ha4, 4'h6 }: pattern = 8'b01100110; 
    { 8'ha4, 4'h7 }: pattern = 8'b01100110; 
    { 8'ha4, 4'h8 }: pattern = 8'b01100110; 
    { 8'ha4, 4'h9 }: pattern = 8'b01100110; 
    { 8'ha4, 4'ha }: pattern = 8'b01100110; 
    { 8'ha4, 4'hb }: pattern = 8'b01100110; 
    { 8'ha4, 4'hc }: pattern = 8'b00000000; 
    { 8'ha4, 4'hd }: pattern = 8'b00000000; 
    { 8'ha4, 4'he }: pattern = 8'b00000000; 
    { 8'ha4, 4'hf }: pattern = 8'b00000000; 

    { 8'ha5, 4'h0 }: pattern = 8'b01110110; 
    { 8'ha5, 4'h1 }: pattern = 8'b11011100; 
    { 8'ha5, 4'h2 }: pattern = 8'b00000000; 
    { 8'ha5, 4'h3 }: pattern = 8'b11000110; 
    { 8'ha5, 4'h4 }: pattern = 8'b11100110; 
    { 8'ha5, 4'h5 }: pattern = 8'b11110110; 
    { 8'ha5, 4'h6 }: pattern = 8'b11111110; 
    { 8'ha5, 4'h7 }: pattern = 8'b11011110; 
    { 8'ha5, 4'h8 }: pattern = 8'b11001110; 
    { 8'ha5, 4'h9 }: pattern = 8'b11000110; 
    { 8'ha5, 4'ha }: pattern = 8'b11000110; 
    { 8'ha5, 4'hb }: pattern = 8'b11000110; 
    { 8'ha5, 4'hc }: pattern = 8'b00000000; 
    { 8'ha5, 4'hd }: pattern = 8'b00000000; 
    { 8'ha5, 4'he }: pattern = 8'b00000000; 
    { 8'ha5, 4'hf }: pattern = 8'b00000000; 

    { 8'ha6, 4'h0 }: pattern = 8'b00000000; 
    { 8'ha6, 4'h1 }: pattern = 8'b00111100; 
    { 8'ha6, 4'h2 }: pattern = 8'b01101100; 
    { 8'ha6, 4'h3 }: pattern = 8'b01101100; 
    { 8'ha6, 4'h4 }: pattern = 8'b00111110; 
    { 8'ha6, 4'h5 }: pattern = 8'b00000000; 
    { 8'ha6, 4'h6 }: pattern = 8'b01111110; 
    { 8'ha6, 4'h7 }: pattern = 8'b00000000; 
    { 8'ha6, 4'h8 }: pattern = 8'b00000000; 
    { 8'ha6, 4'h9 }: pattern = 8'b00000000; 
    { 8'ha6, 4'ha }: pattern = 8'b00000000; 
    { 8'ha6, 4'hb }: pattern = 8'b00000000; 
    { 8'ha6, 4'hc }: pattern = 8'b00000000; 
    { 8'ha6, 4'hd }: pattern = 8'b00000000; 
    { 8'ha6, 4'he }: pattern = 8'b00000000; 
    { 8'ha6, 4'hf }: pattern = 8'b00000000; 

    { 8'ha7, 4'h0 }: pattern = 8'b00000000; 
    { 8'ha7, 4'h1 }: pattern = 8'b00111000; 
    { 8'ha7, 4'h2 }: pattern = 8'b01101100; 
    { 8'ha7, 4'h3 }: pattern = 8'b01101100; 
    { 8'ha7, 4'h4 }: pattern = 8'b00111000; 
    { 8'ha7, 4'h5 }: pattern = 8'b00000000; 
    { 8'ha7, 4'h6 }: pattern = 8'b01111100; 
    { 8'ha7, 4'h7 }: pattern = 8'b00000000; 
    { 8'ha7, 4'h8 }: pattern = 8'b00000000; 
    { 8'ha7, 4'h9 }: pattern = 8'b00000000; 
    { 8'ha7, 4'ha }: pattern = 8'b00000000; 
    { 8'ha7, 4'hb }: pattern = 8'b00000000; 
    { 8'ha7, 4'hc }: pattern = 8'b00000000; 
    { 8'ha7, 4'hd }: pattern = 8'b00000000; 
    { 8'ha7, 4'he }: pattern = 8'b00000000; 
    { 8'ha7, 4'hf }: pattern = 8'b00000000; 

    { 8'ha8, 4'h0 }: pattern = 8'b00000000; 
    { 8'ha8, 4'h1 }: pattern = 8'b00000000; 
    { 8'ha8, 4'h2 }: pattern = 8'b00110000; 
    { 8'ha8, 4'h3 }: pattern = 8'b00110000; 
    { 8'ha8, 4'h4 }: pattern = 8'b00000000; 
    { 8'ha8, 4'h5 }: pattern = 8'b00110000; 
    { 8'ha8, 4'h6 }: pattern = 8'b00110000; 
    { 8'ha8, 4'h7 }: pattern = 8'b01100000; 
    { 8'ha8, 4'h8 }: pattern = 8'b11000000; 
    { 8'ha8, 4'h9 }: pattern = 8'b11000110; 
    { 8'ha8, 4'ha }: pattern = 8'b11000110; 
    { 8'ha8, 4'hb }: pattern = 8'b01111100; 
    { 8'ha8, 4'hc }: pattern = 8'b00000000; 
    { 8'ha8, 4'hd }: pattern = 8'b00000000; 
    { 8'ha8, 4'he }: pattern = 8'b00000000; 
    { 8'ha8, 4'hf }: pattern = 8'b00000000; 

    { 8'ha9, 4'h0 }: pattern = 8'b00000000; 
    { 8'ha9, 4'h1 }: pattern = 8'b00000000; 
    { 8'ha9, 4'h2 }: pattern = 8'b00000000; 
    { 8'ha9, 4'h3 }: pattern = 8'b00000000; 
    { 8'ha9, 4'h4 }: pattern = 8'b00000000; 
    { 8'ha9, 4'h5 }: pattern = 8'b00000000; 
    { 8'ha9, 4'h6 }: pattern = 8'b11111110; 
    { 8'ha9, 4'h7 }: pattern = 8'b11000000; 
    { 8'ha9, 4'h8 }: pattern = 8'b11000000; 
    { 8'ha9, 4'h9 }: pattern = 8'b11000000; 
    { 8'ha9, 4'ha }: pattern = 8'b11000000; 
    { 8'ha9, 4'hb }: pattern = 8'b00000000; 
    { 8'ha9, 4'hc }: pattern = 8'b00000000; 
    { 8'ha9, 4'hd }: pattern = 8'b00000000; 
    { 8'ha9, 4'he }: pattern = 8'b00000000; 
    { 8'ha9, 4'hf }: pattern = 8'b00000000; 

    { 8'haa, 4'h0 }: pattern = 8'b00000000; 
    { 8'haa, 4'h1 }: pattern = 8'b00000000; 
    { 8'haa, 4'h2 }: pattern = 8'b00000000; 
    { 8'haa, 4'h3 }: pattern = 8'b00000000; 
    { 8'haa, 4'h4 }: pattern = 8'b00000000; 
    { 8'haa, 4'h5 }: pattern = 8'b00000000; 
    { 8'haa, 4'h6 }: pattern = 8'b11111110; 
    { 8'haa, 4'h7 }: pattern = 8'b00000110; 
    { 8'haa, 4'h8 }: pattern = 8'b00000110; 
    { 8'haa, 4'h9 }: pattern = 8'b00000110; 
    { 8'haa, 4'ha }: pattern = 8'b00000110; 
    { 8'haa, 4'hb }: pattern = 8'b00000000; 
    { 8'haa, 4'hc }: pattern = 8'b00000000; 
    { 8'haa, 4'hd }: pattern = 8'b00000000; 
    { 8'haa, 4'he }: pattern = 8'b00000000; 
    { 8'haa, 4'hf }: pattern = 8'b00000000; 

    { 8'hab, 4'h0 }: pattern = 8'b00000000; 
    { 8'hab, 4'h1 }: pattern = 8'b11000000; 
    { 8'hab, 4'h2 }: pattern = 8'b11000000; 
    { 8'hab, 4'h3 }: pattern = 8'b11000010; 
    { 8'hab, 4'h4 }: pattern = 8'b11000110; 
    { 8'hab, 4'h5 }: pattern = 8'b11001100; 
    { 8'hab, 4'h6 }: pattern = 8'b00011000; 
    { 8'hab, 4'h7 }: pattern = 8'b00110000; 
    { 8'hab, 4'h8 }: pattern = 8'b01100000; 
    { 8'hab, 4'h9 }: pattern = 8'b11011100; 
    { 8'hab, 4'ha }: pattern = 8'b10000110; 
    { 8'hab, 4'hb }: pattern = 8'b00001100; 
    { 8'hab, 4'hc }: pattern = 8'b00011000; 
    { 8'hab, 4'hd }: pattern = 8'b00111110; 
    { 8'hab, 4'he }: pattern = 8'b00000000; 
    { 8'hab, 4'hf }: pattern = 8'b00000000; 

    { 8'hac, 4'h0 }: pattern = 8'b00000000; 
    { 8'hac, 4'h1 }: pattern = 8'b11000000; 
    { 8'hac, 4'h2 }: pattern = 8'b11000000; 
    { 8'hac, 4'h3 }: pattern = 8'b11000010; 
    { 8'hac, 4'h4 }: pattern = 8'b11000110; 
    { 8'hac, 4'h5 }: pattern = 8'b11001100; 
    { 8'hac, 4'h6 }: pattern = 8'b00011000; 
    { 8'hac, 4'h7 }: pattern = 8'b00110000; 
    { 8'hac, 4'h8 }: pattern = 8'b01100110; 
    { 8'hac, 4'h9 }: pattern = 8'b11001110; 
    { 8'hac, 4'ha }: pattern = 8'b10011110; 
    { 8'hac, 4'hb }: pattern = 8'b00111110; 
    { 8'hac, 4'hc }: pattern = 8'b00000110; 
    { 8'hac, 4'hd }: pattern = 8'b00000110; 
    { 8'hac, 4'he }: pattern = 8'b00000000; 
    { 8'hac, 4'hf }: pattern = 8'b00000000; 

    { 8'had, 4'h0 }: pattern = 8'b00000000; 
    { 8'had, 4'h1 }: pattern = 8'b00000000; 
    { 8'had, 4'h2 }: pattern = 8'b00011000; 
    { 8'had, 4'h3 }: pattern = 8'b00011000; 
    { 8'had, 4'h4 }: pattern = 8'b00000000; 
    { 8'had, 4'h5 }: pattern = 8'b00011000; 
    { 8'had, 4'h6 }: pattern = 8'b00011000; 
    { 8'had, 4'h7 }: pattern = 8'b00011000; 
    { 8'had, 4'h8 }: pattern = 8'b00111100; 
    { 8'had, 4'h9 }: pattern = 8'b00111100; 
    { 8'had, 4'ha }: pattern = 8'b00111100; 
    { 8'had, 4'hb }: pattern = 8'b00011000; 
    { 8'had, 4'hc }: pattern = 8'b00000000; 
    { 8'had, 4'hd }: pattern = 8'b00000000; 
    { 8'had, 4'he }: pattern = 8'b00000000; 
    { 8'had, 4'hf }: pattern = 8'b00000000; 

    { 8'hae, 4'h0 }: pattern = 8'b00000000; 
    { 8'hae, 4'h1 }: pattern = 8'b00000000; 
    { 8'hae, 4'h2 }: pattern = 8'b00000000; 
    { 8'hae, 4'h3 }: pattern = 8'b00000000; 
    { 8'hae, 4'h4 }: pattern = 8'b00000000; 
    { 8'hae, 4'h5 }: pattern = 8'b00110110; 
    { 8'hae, 4'h6 }: pattern = 8'b01101100; 
    { 8'hae, 4'h7 }: pattern = 8'b11011000; 
    { 8'hae, 4'h8 }: pattern = 8'b01101100; 
    { 8'hae, 4'h9 }: pattern = 8'b00110110; 
    { 8'hae, 4'ha }: pattern = 8'b00000000; 
    { 8'hae, 4'hb }: pattern = 8'b00000000; 
    { 8'hae, 4'hc }: pattern = 8'b00000000; 
    { 8'hae, 4'hd }: pattern = 8'b00000000; 
    { 8'hae, 4'he }: pattern = 8'b00000000; 
    { 8'hae, 4'hf }: pattern = 8'b00000000; 

    { 8'haf, 4'h0 }: pattern = 8'b00000000; 
    { 8'haf, 4'h1 }: pattern = 8'b00000000; 
    { 8'haf, 4'h2 }: pattern = 8'b00000000; 
    { 8'haf, 4'h3 }: pattern = 8'b00000000; 
    { 8'haf, 4'h4 }: pattern = 8'b00000000; 
    { 8'haf, 4'h5 }: pattern = 8'b11011000; 
    { 8'haf, 4'h6 }: pattern = 8'b01101100; 
    { 8'haf, 4'h7 }: pattern = 8'b00110110; 
    { 8'haf, 4'h8 }: pattern = 8'b01101100; 
    { 8'haf, 4'h9 }: pattern = 8'b11011000; 
    { 8'haf, 4'ha }: pattern = 8'b00000000; 
    { 8'haf, 4'hb }: pattern = 8'b00000000; 
    { 8'haf, 4'hc }: pattern = 8'b00000000; 
    { 8'haf, 4'hd }: pattern = 8'b00000000; 
    { 8'haf, 4'he }: pattern = 8'b00000000; 
    { 8'haf, 4'hf }: pattern = 8'b00000000; 

    { 8'hb0, 4'h0 }: pattern = 8'b00010001; 
    { 8'hb0, 4'h1 }: pattern = 8'b01000100; 
    { 8'hb0, 4'h2 }: pattern = 8'b00010001; 
    { 8'hb0, 4'h3 }: pattern = 8'b01000100; 
    { 8'hb0, 4'h4 }: pattern = 8'b00010001; 
    { 8'hb0, 4'h5 }: pattern = 8'b01000100; 
    { 8'hb0, 4'h6 }: pattern = 8'b00010001; 
    { 8'hb0, 4'h7 }: pattern = 8'b01000100; 
    { 8'hb0, 4'h8 }: pattern = 8'b00010001; 
    { 8'hb0, 4'h9 }: pattern = 8'b01000100; 
    { 8'hb0, 4'ha }: pattern = 8'b00010001; 
    { 8'hb0, 4'hb }: pattern = 8'b01000100; 
    { 8'hb0, 4'hc }: pattern = 8'b00010001; 
    { 8'hb0, 4'hd }: pattern = 8'b01000100; 
    { 8'hb0, 4'he }: pattern = 8'b00010001; 
    { 8'hb0, 4'hf }: pattern = 8'b01000100; 

    { 8'hb1, 4'h0 }: pattern = 8'b01010101; 
    { 8'hb1, 4'h1 }: pattern = 8'b10101010; 
    { 8'hb1, 4'h2 }: pattern = 8'b01010101; 
    { 8'hb1, 4'h3 }: pattern = 8'b10101010; 
    { 8'hb1, 4'h4 }: pattern = 8'b01010101; 
    { 8'hb1, 4'h5 }: pattern = 8'b10101010; 
    { 8'hb1, 4'h6 }: pattern = 8'b01010101; 
    { 8'hb1, 4'h7 }: pattern = 8'b10101010; 
    { 8'hb1, 4'h8 }: pattern = 8'b01010101; 
    { 8'hb1, 4'h9 }: pattern = 8'b10101010; 
    { 8'hb1, 4'ha }: pattern = 8'b01010101; 
    { 8'hb1, 4'hb }: pattern = 8'b10101010; 
    { 8'hb1, 4'hc }: pattern = 8'b01010101; 
    { 8'hb1, 4'hd }: pattern = 8'b10101010; 
    { 8'hb1, 4'he }: pattern = 8'b01010101; 
    { 8'hb1, 4'hf }: pattern = 8'b10101010; 

    { 8'hb2, 4'h0 }: pattern = 8'b11011101; 
    { 8'hb2, 4'h1 }: pattern = 8'b01110111; 
    { 8'hb2, 4'h2 }: pattern = 8'b11011101; 
    { 8'hb2, 4'h3 }: pattern = 8'b01110111; 
    { 8'hb2, 4'h4 }: pattern = 8'b11011101; 
    { 8'hb2, 4'h5 }: pattern = 8'b01110111; 
    { 8'hb2, 4'h6 }: pattern = 8'b11011101; 
    { 8'hb2, 4'h7 }: pattern = 8'b01110111; 
    { 8'hb2, 4'h8 }: pattern = 8'b11011101; 
    { 8'hb2, 4'h9 }: pattern = 8'b01110111; 
    { 8'hb2, 4'ha }: pattern = 8'b11011101; 
    { 8'hb2, 4'hb }: pattern = 8'b01110111; 
    { 8'hb2, 4'hc }: pattern = 8'b11011101; 
    { 8'hb2, 4'hd }: pattern = 8'b01110111; 
    { 8'hb2, 4'he }: pattern = 8'b11011101; 
    { 8'hb2, 4'hf }: pattern = 8'b01110111; 

    { 8'hb3, 4'h0 }: pattern = 8'b00011000; 
    { 8'hb3, 4'h1 }: pattern = 8'b00011000; 
    { 8'hb3, 4'h2 }: pattern = 8'b00011000; 
    { 8'hb3, 4'h3 }: pattern = 8'b00011000; 
    { 8'hb3, 4'h4 }: pattern = 8'b00011000; 
    { 8'hb3, 4'h5 }: pattern = 8'b00011000; 
    { 8'hb3, 4'h6 }: pattern = 8'b00011000; 
    { 8'hb3, 4'h7 }: pattern = 8'b00011000; 
    { 8'hb3, 4'h8 }: pattern = 8'b00011000; 
    { 8'hb3, 4'h9 }: pattern = 8'b00011000; 
    { 8'hb3, 4'ha }: pattern = 8'b00011000; 
    { 8'hb3, 4'hb }: pattern = 8'b00011000; 
    { 8'hb3, 4'hc }: pattern = 8'b00011000; 
    { 8'hb3, 4'hd }: pattern = 8'b00011000; 
    { 8'hb3, 4'he }: pattern = 8'b00011000; 
    { 8'hb3, 4'hf }: pattern = 8'b00011000; 

    { 8'hb4, 4'h0 }: pattern = 8'b00011000; 
    { 8'hb4, 4'h1 }: pattern = 8'b00011000; 
    { 8'hb4, 4'h2 }: pattern = 8'b00011000; 
    { 8'hb4, 4'h3 }: pattern = 8'b00011000; 
    { 8'hb4, 4'h4 }: pattern = 8'b00011000; 
    { 8'hb4, 4'h5 }: pattern = 8'b00011000; 
    { 8'hb4, 4'h6 }: pattern = 8'b00011000; 
    { 8'hb4, 4'h7 }: pattern = 8'b11111000; 
    { 8'hb4, 4'h8 }: pattern = 8'b00011000; 
    { 8'hb4, 4'h9 }: pattern = 8'b00011000; 
    { 8'hb4, 4'ha }: pattern = 8'b00011000; 
    { 8'hb4, 4'hb }: pattern = 8'b00011000; 
    { 8'hb4, 4'hc }: pattern = 8'b00011000; 
    { 8'hb4, 4'hd }: pattern = 8'b00011000; 
    { 8'hb4, 4'he }: pattern = 8'b00011000; 
    { 8'hb4, 4'hf }: pattern = 8'b00011000; 

    { 8'hb5, 4'h0 }: pattern = 8'b00011000; 
    { 8'hb5, 4'h1 }: pattern = 8'b00011000; 
    { 8'hb5, 4'h2 }: pattern = 8'b00011000; 
    { 8'hb5, 4'h3 }: pattern = 8'b00011000; 
    { 8'hb5, 4'h4 }: pattern = 8'b00011000; 
    { 8'hb5, 4'h5 }: pattern = 8'b11111000; 
    { 8'hb5, 4'h6 }: pattern = 8'b00011000; 
    { 8'hb5, 4'h7 }: pattern = 8'b11111000; 
    { 8'hb5, 4'h8 }: pattern = 8'b00011000; 
    { 8'hb5, 4'h9 }: pattern = 8'b00011000; 
    { 8'hb5, 4'ha }: pattern = 8'b00011000; 
    { 8'hb5, 4'hb }: pattern = 8'b00011000; 
    { 8'hb5, 4'hc }: pattern = 8'b00011000; 
    { 8'hb5, 4'hd }: pattern = 8'b00011000; 
    { 8'hb5, 4'he }: pattern = 8'b00011000; 
    { 8'hb5, 4'hf }: pattern = 8'b00011000; 

    { 8'hb6, 4'h0 }: pattern = 8'b00110110; 
    { 8'hb6, 4'h1 }: pattern = 8'b00110110; 
    { 8'hb6, 4'h2 }: pattern = 8'b00110110; 
    { 8'hb6, 4'h3 }: pattern = 8'b00110110; 
    { 8'hb6, 4'h4 }: pattern = 8'b00110110; 
    { 8'hb6, 4'h5 }: pattern = 8'b00110110; 
    { 8'hb6, 4'h6 }: pattern = 8'b00110110; 
    { 8'hb6, 4'h7 }: pattern = 8'b11110110; 
    { 8'hb6, 4'h8 }: pattern = 8'b00110110; 
    { 8'hb6, 4'h9 }: pattern = 8'b00110110; 
    { 8'hb6, 4'ha }: pattern = 8'b00110110; 
    { 8'hb6, 4'hb }: pattern = 8'b00110110; 
    { 8'hb6, 4'hc }: pattern = 8'b00110110; 
    { 8'hb6, 4'hd }: pattern = 8'b00110110; 
    { 8'hb6, 4'he }: pattern = 8'b00110110; 
    { 8'hb6, 4'hf }: pattern = 8'b00110110; 

    { 8'hb7, 4'h0 }: pattern = 8'b00000000; 
    { 8'hb7, 4'h1 }: pattern = 8'b00000000; 
    { 8'hb7, 4'h2 }: pattern = 8'b00000000; 
    { 8'hb7, 4'h3 }: pattern = 8'b00000000; 
    { 8'hb7, 4'h4 }: pattern = 8'b00000000; 
    { 8'hb7, 4'h5 }: pattern = 8'b00000000; 
    { 8'hb7, 4'h6 }: pattern = 8'b00000000; 
    { 8'hb7, 4'h7 }: pattern = 8'b11111110; 
    { 8'hb7, 4'h8 }: pattern = 8'b00110110; 
    { 8'hb7, 4'h9 }: pattern = 8'b00110110; 
    { 8'hb7, 4'ha }: pattern = 8'b00110110; 
    { 8'hb7, 4'hb }: pattern = 8'b00110110; 
    { 8'hb7, 4'hc }: pattern = 8'b00110110; 
    { 8'hb7, 4'hd }: pattern = 8'b00110110; 
    { 8'hb7, 4'he }: pattern = 8'b00110110; 
    { 8'hb7, 4'hf }: pattern = 8'b00110110; 

    { 8'hb8, 4'h0 }: pattern = 8'b00000000; 
    { 8'hb8, 4'h1 }: pattern = 8'b00000000; 
    { 8'hb8, 4'h2 }: pattern = 8'b00000000; 
    { 8'hb8, 4'h3 }: pattern = 8'b00000000; 
    { 8'hb8, 4'h4 }: pattern = 8'b00000000; 
    { 8'hb8, 4'h5 }: pattern = 8'b11111000; 
    { 8'hb8, 4'h6 }: pattern = 8'b00011000; 
    { 8'hb8, 4'h7 }: pattern = 8'b11111000; 
    { 8'hb8, 4'h8 }: pattern = 8'b00011000; 
    { 8'hb8, 4'h9 }: pattern = 8'b00011000; 
    { 8'hb8, 4'ha }: pattern = 8'b00011000; 
    { 8'hb8, 4'hb }: pattern = 8'b00011000; 
    { 8'hb8, 4'hc }: pattern = 8'b00011000; 
    { 8'hb8, 4'hd }: pattern = 8'b00011000; 
    { 8'hb8, 4'he }: pattern = 8'b00011000; 
    { 8'hb8, 4'hf }: pattern = 8'b00011000; 

    { 8'hb9, 4'h0 }: pattern = 8'b00110110; 
    { 8'hb9, 4'h1 }: pattern = 8'b00110110; 
    { 8'hb9, 4'h2 }: pattern = 8'b00110110; 
    { 8'hb9, 4'h3 }: pattern = 8'b00110110; 
    { 8'hb9, 4'h4 }: pattern = 8'b00110110; 
    { 8'hb9, 4'h5 }: pattern = 8'b11110110; 
    { 8'hb9, 4'h6 }: pattern = 8'b00000110; 
    { 8'hb9, 4'h7 }: pattern = 8'b11110110; 
    { 8'hb9, 4'h8 }: pattern = 8'b00110110; 
    { 8'hb9, 4'h9 }: pattern = 8'b00110110; 
    { 8'hb9, 4'ha }: pattern = 8'b00110110; 
    { 8'hb9, 4'hb }: pattern = 8'b00110110; 
    { 8'hb9, 4'hc }: pattern = 8'b00110110; 
    { 8'hb9, 4'hd }: pattern = 8'b00110110; 
    { 8'hb9, 4'he }: pattern = 8'b00110110; 
    { 8'hb9, 4'hf }: pattern = 8'b00110110; 

    { 8'hba, 4'h0 }: pattern = 8'b00110110; 
    { 8'hba, 4'h1 }: pattern = 8'b00110110; 
    { 8'hba, 4'h2 }: pattern = 8'b00110110; 
    { 8'hba, 4'h3 }: pattern = 8'b00110110; 
    { 8'hba, 4'h4 }: pattern = 8'b00110110; 
    { 8'hba, 4'h5 }: pattern = 8'b00110110; 
    { 8'hba, 4'h6 }: pattern = 8'b00110110; 
    { 8'hba, 4'h7 }: pattern = 8'b00110110; 
    { 8'hba, 4'h8 }: pattern = 8'b00110110; 
    { 8'hba, 4'h9 }: pattern = 8'b00110110; 
    { 8'hba, 4'ha }: pattern = 8'b00110110; 
    { 8'hba, 4'hb }: pattern = 8'b00110110; 
    { 8'hba, 4'hc }: pattern = 8'b00110110; 
    { 8'hba, 4'hd }: pattern = 8'b00110110; 
    { 8'hba, 4'he }: pattern = 8'b00110110; 
    { 8'hba, 4'hf }: pattern = 8'b00110110; 

    { 8'hbb, 4'h0 }: pattern = 8'b00000000; 
    { 8'hbb, 4'h1 }: pattern = 8'b00000000; 
    { 8'hbb, 4'h2 }: pattern = 8'b00000000; 
    { 8'hbb, 4'h3 }: pattern = 8'b00000000; 
    { 8'hbb, 4'h4 }: pattern = 8'b00000000; 
    { 8'hbb, 4'h5 }: pattern = 8'b11111110; 
    { 8'hbb, 4'h6 }: pattern = 8'b00000110; 
    { 8'hbb, 4'h7 }: pattern = 8'b11110110; 
    { 8'hbb, 4'h8 }: pattern = 8'b00110110; 
    { 8'hbb, 4'h9 }: pattern = 8'b00110110; 
    { 8'hbb, 4'ha }: pattern = 8'b00110110; 
    { 8'hbb, 4'hb }: pattern = 8'b00110110; 
    { 8'hbb, 4'hc }: pattern = 8'b00110110; 
    { 8'hbb, 4'hd }: pattern = 8'b00110110; 
    { 8'hbb, 4'he }: pattern = 8'b00110110; 
    { 8'hbb, 4'hf }: pattern = 8'b00110110; 

    { 8'hbc, 4'h0 }: pattern = 8'b00110110; 
    { 8'hbc, 4'h1 }: pattern = 8'b00110110; 
    { 8'hbc, 4'h2 }: pattern = 8'b00110110; 
    { 8'hbc, 4'h3 }: pattern = 8'b00110110; 
    { 8'hbc, 4'h4 }: pattern = 8'b00110110; 
    { 8'hbc, 4'h5 }: pattern = 8'b11110110; 
    { 8'hbc, 4'h6 }: pattern = 8'b00000110; 
    { 8'hbc, 4'h7 }: pattern = 8'b11111110; 
    { 8'hbc, 4'h8 }: pattern = 8'b00000000; 
    { 8'hbc, 4'h9 }: pattern = 8'b00000000; 
    { 8'hbc, 4'ha }: pattern = 8'b00000000; 
    { 8'hbc, 4'hb }: pattern = 8'b00000000; 
    { 8'hbc, 4'hc }: pattern = 8'b00000000; 
    { 8'hbc, 4'hd }: pattern = 8'b00000000; 
    { 8'hbc, 4'he }: pattern = 8'b00000000; 
    { 8'hbc, 4'hf }: pattern = 8'b00000000; 

    { 8'hbd, 4'h0 }: pattern = 8'b00110110; 
    { 8'hbd, 4'h1 }: pattern = 8'b00110110; 
    { 8'hbd, 4'h2 }: pattern = 8'b00110110; 
    { 8'hbd, 4'h3 }: pattern = 8'b00110110; 
    { 8'hbd, 4'h4 }: pattern = 8'b00110110; 
    { 8'hbd, 4'h5 }: pattern = 8'b00110110; 
    { 8'hbd, 4'h6 }: pattern = 8'b00110110; 
    { 8'hbd, 4'h7 }: pattern = 8'b11111110; 
    { 8'hbd, 4'h8 }: pattern = 8'b00000000; 
    { 8'hbd, 4'h9 }: pattern = 8'b00000000; 
    { 8'hbd, 4'ha }: pattern = 8'b00000000; 
    { 8'hbd, 4'hb }: pattern = 8'b00000000; 
    { 8'hbd, 4'hc }: pattern = 8'b00000000; 
    { 8'hbd, 4'hd }: pattern = 8'b00000000; 
    { 8'hbd, 4'he }: pattern = 8'b00000000; 
    { 8'hbd, 4'hf }: pattern = 8'b00000000; 

    { 8'hbe, 4'h0 }: pattern = 8'b00011000; 
    { 8'hbe, 4'h1 }: pattern = 8'b00011000; 
    { 8'hbe, 4'h2 }: pattern = 8'b00011000; 
    { 8'hbe, 4'h3 }: pattern = 8'b00011000; 
    { 8'hbe, 4'h4 }: pattern = 8'b00011000; 
    { 8'hbe, 4'h5 }: pattern = 8'b11111000; 
    { 8'hbe, 4'h6 }: pattern = 8'b00011000; 
    { 8'hbe, 4'h7 }: pattern = 8'b11111000; 
    { 8'hbe, 4'h8 }: pattern = 8'b00000000; 
    { 8'hbe, 4'h9 }: pattern = 8'b00000000; 
    { 8'hbe, 4'ha }: pattern = 8'b00000000; 
    { 8'hbe, 4'hb }: pattern = 8'b00000000; 
    { 8'hbe, 4'hc }: pattern = 8'b00000000; 
    { 8'hbe, 4'hd }: pattern = 8'b00000000; 
    { 8'hbe, 4'he }: pattern = 8'b00000000; 
    { 8'hbe, 4'hf }: pattern = 8'b00000000; 

    { 8'hbf, 4'h0 }: pattern = 8'b00000000; 
    { 8'hbf, 4'h1 }: pattern = 8'b00000000; 
    { 8'hbf, 4'h2 }: pattern = 8'b00000000; 
    { 8'hbf, 4'h3 }: pattern = 8'b00000000; 
    { 8'hbf, 4'h4 }: pattern = 8'b00000000; 
    { 8'hbf, 4'h5 }: pattern = 8'b00000000; 
    { 8'hbf, 4'h6 }: pattern = 8'b00000000; 
    { 8'hbf, 4'h7 }: pattern = 8'b11111000; 
    { 8'hbf, 4'h8 }: pattern = 8'b00011000; 
    { 8'hbf, 4'h9 }: pattern = 8'b00011000; 
    { 8'hbf, 4'ha }: pattern = 8'b00011000; 
    { 8'hbf, 4'hb }: pattern = 8'b00011000; 
    { 8'hbf, 4'hc }: pattern = 8'b00011000; 
    { 8'hbf, 4'hd }: pattern = 8'b00011000; 
    { 8'hbf, 4'he }: pattern = 8'b00011000; 
    { 8'hbf, 4'hf }: pattern = 8'b00011000; 

    { 8'hc0, 4'h0 }: pattern = 8'b00011000; 
    { 8'hc0, 4'h1 }: pattern = 8'b00011000; 
    { 8'hc0, 4'h2 }: pattern = 8'b00011000; 
    { 8'hc0, 4'h3 }: pattern = 8'b00011000; 
    { 8'hc0, 4'h4 }: pattern = 8'b00011000; 
    { 8'hc0, 4'h5 }: pattern = 8'b00011000; 
    { 8'hc0, 4'h6 }: pattern = 8'b00011000; 
    { 8'hc0, 4'h7 }: pattern = 8'b00011111; 
    { 8'hc0, 4'h8 }: pattern = 8'b00000000; 
    { 8'hc0, 4'h9 }: pattern = 8'b00000000; 
    { 8'hc0, 4'ha }: pattern = 8'b00000000; 
    { 8'hc0, 4'hb }: pattern = 8'b00000000; 
    { 8'hc0, 4'hc }: pattern = 8'b00000000; 
    { 8'hc0, 4'hd }: pattern = 8'b00000000; 
    { 8'hc0, 4'he }: pattern = 8'b00000000; 
    { 8'hc0, 4'hf }: pattern = 8'b00000000; 

    { 8'hc1, 4'h0 }: pattern = 8'b00011000; 
    { 8'hc1, 4'h1 }: pattern = 8'b00011000; 
    { 8'hc1, 4'h2 }: pattern = 8'b00011000; 
    { 8'hc1, 4'h3 }: pattern = 8'b00011000; 
    { 8'hc1, 4'h4 }: pattern = 8'b00011000; 
    { 8'hc1, 4'h5 }: pattern = 8'b00011000; 
    { 8'hc1, 4'h6 }: pattern = 8'b00011000; 
    { 8'hc1, 4'h7 }: pattern = 8'b11111111; 
    { 8'hc1, 4'h8 }: pattern = 8'b00000000; 
    { 8'hc1, 4'h9 }: pattern = 8'b00000000; 
    { 8'hc1, 4'ha }: pattern = 8'b00000000; 
    { 8'hc1, 4'hb }: pattern = 8'b00000000; 
    { 8'hc1, 4'hc }: pattern = 8'b00000000; 
    { 8'hc1, 4'hd }: pattern = 8'b00000000; 
    { 8'hc1, 4'he }: pattern = 8'b00000000; 
    { 8'hc1, 4'hf }: pattern = 8'b00000000; 

    { 8'hc2, 4'h0 }: pattern = 8'b00000000; 
    { 8'hc2, 4'h1 }: pattern = 8'b00000000; 
    { 8'hc2, 4'h2 }: pattern = 8'b00000000; 
    { 8'hc2, 4'h3 }: pattern = 8'b00000000; 
    { 8'hc2, 4'h4 }: pattern = 8'b00000000; 
    { 8'hc2, 4'h5 }: pattern = 8'b00000000; 
    { 8'hc2, 4'h6 }: pattern = 8'b00000000; 
    { 8'hc2, 4'h7 }: pattern = 8'b11111111; 
    { 8'hc2, 4'h8 }: pattern = 8'b00011000; 
    { 8'hc2, 4'h9 }: pattern = 8'b00011000; 
    { 8'hc2, 4'ha }: pattern = 8'b00011000; 
    { 8'hc2, 4'hb }: pattern = 8'b00011000; 
    { 8'hc2, 4'hc }: pattern = 8'b00011000; 
    { 8'hc2, 4'hd }: pattern = 8'b00011000; 
    { 8'hc2, 4'he }: pattern = 8'b00011000; 
    { 8'hc2, 4'hf }: pattern = 8'b00011000; 

    { 8'hc3, 4'h0 }: pattern = 8'b00011000; 
    { 8'hc3, 4'h1 }: pattern = 8'b00011000; 
    { 8'hc3, 4'h2 }: pattern = 8'b00011000; 
    { 8'hc3, 4'h3 }: pattern = 8'b00011000; 
    { 8'hc3, 4'h4 }: pattern = 8'b00011000; 
    { 8'hc3, 4'h5 }: pattern = 8'b00011000; 
    { 8'hc3, 4'h6 }: pattern = 8'b00011000; 
    { 8'hc3, 4'h7 }: pattern = 8'b00011111; 
    { 8'hc3, 4'h8 }: pattern = 8'b00011000; 
    { 8'hc3, 4'h9 }: pattern = 8'b00011000; 
    { 8'hc3, 4'ha }: pattern = 8'b00011000; 
    { 8'hc3, 4'hb }: pattern = 8'b00011000; 
    { 8'hc3, 4'hc }: pattern = 8'b00011000; 
    { 8'hc3, 4'hd }: pattern = 8'b00011000; 
    { 8'hc3, 4'he }: pattern = 8'b00011000; 
    { 8'hc3, 4'hf }: pattern = 8'b00011000; 

    { 8'hc4, 4'h0 }: pattern = 8'b00000000; 
    { 8'hc4, 4'h1 }: pattern = 8'b00000000; 
    { 8'hc4, 4'h2 }: pattern = 8'b00000000; 
    { 8'hc4, 4'h3 }: pattern = 8'b00000000; 
    { 8'hc4, 4'h4 }: pattern = 8'b00000000; 
    { 8'hc4, 4'h5 }: pattern = 8'b00000000; 
    { 8'hc4, 4'h6 }: pattern = 8'b00000000; 
    { 8'hc4, 4'h7 }: pattern = 8'b11111111; 
    { 8'hc4, 4'h8 }: pattern = 8'b00000000; 
    { 8'hc4, 4'h9 }: pattern = 8'b00000000; 
    { 8'hc4, 4'ha }: pattern = 8'b00000000; 
    { 8'hc4, 4'hb }: pattern = 8'b00000000; 
    { 8'hc4, 4'hc }: pattern = 8'b00000000; 
    { 8'hc4, 4'hd }: pattern = 8'b00000000; 
    { 8'hc4, 4'he }: pattern = 8'b00000000; 
    { 8'hc4, 4'hf }: pattern = 8'b00000000; 

    { 8'hc5, 4'h0 }: pattern = 8'b00011000; 
    { 8'hc5, 4'h1 }: pattern = 8'b00011000; 
    { 8'hc5, 4'h2 }: pattern = 8'b00011000; 
    { 8'hc5, 4'h3 }: pattern = 8'b00011000; 
    { 8'hc5, 4'h4 }: pattern = 8'b00011000; 
    { 8'hc5, 4'h5 }: pattern = 8'b00011000; 
    { 8'hc5, 4'h6 }: pattern = 8'b00011000; 
    { 8'hc5, 4'h7 }: pattern = 8'b11111111; 
    { 8'hc5, 4'h8 }: pattern = 8'b00011000; 
    { 8'hc5, 4'h9 }: pattern = 8'b00011000; 
    { 8'hc5, 4'ha }: pattern = 8'b00011000; 
    { 8'hc5, 4'hb }: pattern = 8'b00011000; 
    { 8'hc5, 4'hc }: pattern = 8'b00011000; 
    { 8'hc5, 4'hd }: pattern = 8'b00011000; 
    { 8'hc5, 4'he }: pattern = 8'b00011000; 
    { 8'hc5, 4'hf }: pattern = 8'b00011000; 

    { 8'hc6, 4'h0 }: pattern = 8'b00011000; 
    { 8'hc6, 4'h1 }: pattern = 8'b00011000; 
    { 8'hc6, 4'h2 }: pattern = 8'b00011000; 
    { 8'hc6, 4'h3 }: pattern = 8'b00011000; 
    { 8'hc6, 4'h4 }: pattern = 8'b00011000; 
    { 8'hc6, 4'h5 }: pattern = 8'b00011111; 
    { 8'hc6, 4'h6 }: pattern = 8'b00011000; 
    { 8'hc6, 4'h7 }: pattern = 8'b00011111; 
    { 8'hc6, 4'h8 }: pattern = 8'b00011000; 
    { 8'hc6, 4'h9 }: pattern = 8'b00011000; 
    { 8'hc6, 4'ha }: pattern = 8'b00011000; 
    { 8'hc6, 4'hb }: pattern = 8'b00011000; 
    { 8'hc6, 4'hc }: pattern = 8'b00011000; 
    { 8'hc6, 4'hd }: pattern = 8'b00011000; 
    { 8'hc6, 4'he }: pattern = 8'b00011000; 
    { 8'hc6, 4'hf }: pattern = 8'b00011000; 

    { 8'hc7, 4'h0 }: pattern = 8'b00110110; 
    { 8'hc7, 4'h1 }: pattern = 8'b00110110; 
    { 8'hc7, 4'h2 }: pattern = 8'b00110110; 
    { 8'hc7, 4'h3 }: pattern = 8'b00110110; 
    { 8'hc7, 4'h4 }: pattern = 8'b00110110; 
    { 8'hc7, 4'h5 }: pattern = 8'b00110110; 
    { 8'hc7, 4'h6 }: pattern = 8'b00110110; 
    { 8'hc7, 4'h7 }: pattern = 8'b00110111; 
    { 8'hc7, 4'h8 }: pattern = 8'b00110110; 
    { 8'hc7, 4'h9 }: pattern = 8'b00110110; 
    { 8'hc7, 4'ha }: pattern = 8'b00110110; 
    { 8'hc7, 4'hb }: pattern = 8'b00110110; 
    { 8'hc7, 4'hc }: pattern = 8'b00110110; 
    { 8'hc7, 4'hd }: pattern = 8'b00110110; 
    { 8'hc7, 4'he }: pattern = 8'b00110110; 
    { 8'hc7, 4'hf }: pattern = 8'b00110110; 

    { 8'hc8, 4'h0 }: pattern = 8'b00110110; 
    { 8'hc8, 4'h1 }: pattern = 8'b00110110; 
    { 8'hc8, 4'h2 }: pattern = 8'b00110110; 
    { 8'hc8, 4'h3 }: pattern = 8'b00110110; 
    { 8'hc8, 4'h4 }: pattern = 8'b00110110; 
    { 8'hc8, 4'h5 }: pattern = 8'b00110111; 
    { 8'hc8, 4'h6 }: pattern = 8'b00110000; 
    { 8'hc8, 4'h7 }: pattern = 8'b00111111; 
    { 8'hc8, 4'h8 }: pattern = 8'b00000000; 
    { 8'hc8, 4'h9 }: pattern = 8'b00000000; 
    { 8'hc8, 4'ha }: pattern = 8'b00000000; 
    { 8'hc8, 4'hb }: pattern = 8'b00000000; 
    { 8'hc8, 4'hc }: pattern = 8'b00000000; 
    { 8'hc8, 4'hd }: pattern = 8'b00000000; 
    { 8'hc8, 4'he }: pattern = 8'b00000000; 
    { 8'hc8, 4'hf }: pattern = 8'b00000000; 

    { 8'hc9, 4'h0 }: pattern = 8'b00000000; 
    { 8'hc9, 4'h1 }: pattern = 8'b00000000; 
    { 8'hc9, 4'h2 }: pattern = 8'b00000000; 
    { 8'hc9, 4'h3 }: pattern = 8'b00000000; 
    { 8'hc9, 4'h4 }: pattern = 8'b00000000; 
    { 8'hc9, 4'h5 }: pattern = 8'b00111111; 
    { 8'hc9, 4'h6 }: pattern = 8'b00110000; 
    { 8'hc9, 4'h7 }: pattern = 8'b00110111; 
    { 8'hc9, 4'h8 }: pattern = 8'b00110110; 
    { 8'hc9, 4'h9 }: pattern = 8'b00110110; 
    { 8'hc9, 4'ha }: pattern = 8'b00110110; 
    { 8'hc9, 4'hb }: pattern = 8'b00110110; 
    { 8'hc9, 4'hc }: pattern = 8'b00110110; 
    { 8'hc9, 4'hd }: pattern = 8'b00110110; 
    { 8'hc9, 4'he }: pattern = 8'b00110110; 
    { 8'hc9, 4'hf }: pattern = 8'b00110110; 

    { 8'hca, 4'h0 }: pattern = 8'b00110110; 
    { 8'hca, 4'h1 }: pattern = 8'b00110110; 
    { 8'hca, 4'h2 }: pattern = 8'b00110110; 
    { 8'hca, 4'h3 }: pattern = 8'b00110110; 
    { 8'hca, 4'h4 }: pattern = 8'b00110110; 
    { 8'hca, 4'h5 }: pattern = 8'b11110111; 
    { 8'hca, 4'h6 }: pattern = 8'b00000000; 
    { 8'hca, 4'h7 }: pattern = 8'b11111111; 
    { 8'hca, 4'h8 }: pattern = 8'b00000000; 
    { 8'hca, 4'h9 }: pattern = 8'b00000000; 
    { 8'hca, 4'ha }: pattern = 8'b00000000; 
    { 8'hca, 4'hb }: pattern = 8'b00000000; 
    { 8'hca, 4'hc }: pattern = 8'b00000000; 
    { 8'hca, 4'hd }: pattern = 8'b00000000; 
    { 8'hca, 4'he }: pattern = 8'b00000000; 
    { 8'hca, 4'hf }: pattern = 8'b00000000; 

    { 8'hcb, 4'h0 }: pattern = 8'b00000000; 
    { 8'hcb, 4'h1 }: pattern = 8'b00000000; 
    { 8'hcb, 4'h2 }: pattern = 8'b00000000; 
    { 8'hcb, 4'h3 }: pattern = 8'b00000000; 
    { 8'hcb, 4'h4 }: pattern = 8'b00000000; 
    { 8'hcb, 4'h5 }: pattern = 8'b11111111; 
    { 8'hcb, 4'h6 }: pattern = 8'b00000000; 
    { 8'hcb, 4'h7 }: pattern = 8'b11110111; 
    { 8'hcb, 4'h8 }: pattern = 8'b00110110; 
    { 8'hcb, 4'h9 }: pattern = 8'b00110110; 
    { 8'hcb, 4'ha }: pattern = 8'b00110110; 
    { 8'hcb, 4'hb }: pattern = 8'b00110110; 
    { 8'hcb, 4'hc }: pattern = 8'b00110110; 
    { 8'hcb, 4'hd }: pattern = 8'b00110110; 
    { 8'hcb, 4'he }: pattern = 8'b00110110; 
    { 8'hcb, 4'hf }: pattern = 8'b00110110; 

    { 8'hcc, 4'h0 }: pattern = 8'b00110110; 
    { 8'hcc, 4'h1 }: pattern = 8'b00110110; 
    { 8'hcc, 4'h2 }: pattern = 8'b00110110; 
    { 8'hcc, 4'h3 }: pattern = 8'b00110110; 
    { 8'hcc, 4'h4 }: pattern = 8'b00110110; 
    { 8'hcc, 4'h5 }: pattern = 8'b00110111; 
    { 8'hcc, 4'h6 }: pattern = 8'b00110000; 
    { 8'hcc, 4'h7 }: pattern = 8'b00110111; 
    { 8'hcc, 4'h8 }: pattern = 8'b00110110; 
    { 8'hcc, 4'h9 }: pattern = 8'b00110110; 
    { 8'hcc, 4'ha }: pattern = 8'b00110110; 
    { 8'hcc, 4'hb }: pattern = 8'b00110110; 
    { 8'hcc, 4'hc }: pattern = 8'b00110110; 
    { 8'hcc, 4'hd }: pattern = 8'b00110110; 
    { 8'hcc, 4'he }: pattern = 8'b00110110; 
    { 8'hcc, 4'hf }: pattern = 8'b00110110; 

    { 8'hcd, 4'h0 }: pattern = 8'b00000000; 
    { 8'hcd, 4'h1 }: pattern = 8'b00000000; 
    { 8'hcd, 4'h2 }: pattern = 8'b00000000; 
    { 8'hcd, 4'h3 }: pattern = 8'b00000000; 
    { 8'hcd, 4'h4 }: pattern = 8'b00000000; 
    { 8'hcd, 4'h5 }: pattern = 8'b11111111; 
    { 8'hcd, 4'h6 }: pattern = 8'b00000000; 
    { 8'hcd, 4'h7 }: pattern = 8'b11111111; 
    { 8'hcd, 4'h8 }: pattern = 8'b00000000; 
    { 8'hcd, 4'h9 }: pattern = 8'b00000000; 
    { 8'hcd, 4'ha }: pattern = 8'b00000000; 
    { 8'hcd, 4'hb }: pattern = 8'b00000000; 
    { 8'hcd, 4'hc }: pattern = 8'b00000000; 
    { 8'hcd, 4'hd }: pattern = 8'b00000000; 
    { 8'hcd, 4'he }: pattern = 8'b00000000; 
    { 8'hcd, 4'hf }: pattern = 8'b00000000; 

    { 8'hce, 4'h0 }: pattern = 8'b00110110; 
    { 8'hce, 4'h1 }: pattern = 8'b00110110; 
    { 8'hce, 4'h2 }: pattern = 8'b00110110; 
    { 8'hce, 4'h3 }: pattern = 8'b00110110; 
    { 8'hce, 4'h4 }: pattern = 8'b00110110; 
    { 8'hce, 4'h5 }: pattern = 8'b11110111; 
    { 8'hce, 4'h6 }: pattern = 8'b00000000; 
    { 8'hce, 4'h7 }: pattern = 8'b11110111; 
    { 8'hce, 4'h8 }: pattern = 8'b00110110; 
    { 8'hce, 4'h9 }: pattern = 8'b00110110; 
    { 8'hce, 4'ha }: pattern = 8'b00110110; 
    { 8'hce, 4'hb }: pattern = 8'b00110110; 
    { 8'hce, 4'hc }: pattern = 8'b00110110; 
    { 8'hce, 4'hd }: pattern = 8'b00110110; 
    { 8'hce, 4'he }: pattern = 8'b00110110; 
    { 8'hce, 4'hf }: pattern = 8'b00110110; 

    { 8'hcf, 4'h0 }: pattern = 8'b00011000; 
    { 8'hcf, 4'h1 }: pattern = 8'b00011000; 
    { 8'hcf, 4'h2 }: pattern = 8'b00011000; 
    { 8'hcf, 4'h3 }: pattern = 8'b00011000; 
    { 8'hcf, 4'h4 }: pattern = 8'b00011000; 
    { 8'hcf, 4'h5 }: pattern = 8'b11111111; 
    { 8'hcf, 4'h6 }: pattern = 8'b00000000; 
    { 8'hcf, 4'h7 }: pattern = 8'b11111111; 
    { 8'hcf, 4'h8 }: pattern = 8'b00000000; 
    { 8'hcf, 4'h9 }: pattern = 8'b00000000; 
    { 8'hcf, 4'ha }: pattern = 8'b00000000; 
    { 8'hcf, 4'hb }: pattern = 8'b00000000; 
    { 8'hcf, 4'hc }: pattern = 8'b00000000; 
    { 8'hcf, 4'hd }: pattern = 8'b00000000; 
    { 8'hcf, 4'he }: pattern = 8'b00000000; 
    { 8'hcf, 4'hf }: pattern = 8'b00000000; 

    { 8'hd0, 4'h0 }: pattern = 8'b00110110; 
    { 8'hd0, 4'h1 }: pattern = 8'b00110110; 
    { 8'hd0, 4'h2 }: pattern = 8'b00110110; 
    { 8'hd0, 4'h3 }: pattern = 8'b00110110; 
    { 8'hd0, 4'h4 }: pattern = 8'b00110110; 
    { 8'hd0, 4'h5 }: pattern = 8'b00110110; 
    { 8'hd0, 4'h6 }: pattern = 8'b00110110; 
    { 8'hd0, 4'h7 }: pattern = 8'b11111111; 
    { 8'hd0, 4'h8 }: pattern = 8'b00000000; 
    { 8'hd0, 4'h9 }: pattern = 8'b00000000; 
    { 8'hd0, 4'ha }: pattern = 8'b00000000; 
    { 8'hd0, 4'hb }: pattern = 8'b00000000; 
    { 8'hd0, 4'hc }: pattern = 8'b00000000; 
    { 8'hd0, 4'hd }: pattern = 8'b00000000; 
    { 8'hd0, 4'he }: pattern = 8'b00000000; 
    { 8'hd0, 4'hf }: pattern = 8'b00000000; 

    { 8'hd1, 4'h0 }: pattern = 8'b00000000; 
    { 8'hd1, 4'h1 }: pattern = 8'b00000000; 
    { 8'hd1, 4'h2 }: pattern = 8'b00000000; 
    { 8'hd1, 4'h3 }: pattern = 8'b00000000; 
    { 8'hd1, 4'h4 }: pattern = 8'b00000000; 
    { 8'hd1, 4'h5 }: pattern = 8'b11111111; 
    { 8'hd1, 4'h6 }: pattern = 8'b00000000; 
    { 8'hd1, 4'h7 }: pattern = 8'b11111111; 
    { 8'hd1, 4'h8 }: pattern = 8'b00011000; 
    { 8'hd1, 4'h9 }: pattern = 8'b00011000; 
    { 8'hd1, 4'ha }: pattern = 8'b00011000; 
    { 8'hd1, 4'hb }: pattern = 8'b00011000; 
    { 8'hd1, 4'hc }: pattern = 8'b00011000; 
    { 8'hd1, 4'hd }: pattern = 8'b00011000; 
    { 8'hd1, 4'he }: pattern = 8'b00011000; 
    { 8'hd1, 4'hf }: pattern = 8'b00011000; 

    { 8'hd2, 4'h0 }: pattern = 8'b00000000; 
    { 8'hd2, 4'h1 }: pattern = 8'b00000000; 
    { 8'hd2, 4'h2 }: pattern = 8'b00000000; 
    { 8'hd2, 4'h3 }: pattern = 8'b00000000; 
    { 8'hd2, 4'h4 }: pattern = 8'b00000000; 
    { 8'hd2, 4'h5 }: pattern = 8'b00000000; 
    { 8'hd2, 4'h6 }: pattern = 8'b00000000; 
    { 8'hd2, 4'h7 }: pattern = 8'b11111111; 
    { 8'hd2, 4'h8 }: pattern = 8'b00110110; 
    { 8'hd2, 4'h9 }: pattern = 8'b00110110; 
    { 8'hd2, 4'ha }: pattern = 8'b00110110; 
    { 8'hd2, 4'hb }: pattern = 8'b00110110; 
    { 8'hd2, 4'hc }: pattern = 8'b00110110; 
    { 8'hd2, 4'hd }: pattern = 8'b00110110; 
    { 8'hd2, 4'he }: pattern = 8'b00110110; 
    { 8'hd2, 4'hf }: pattern = 8'b00110110; 

    { 8'hd3, 4'h0 }: pattern = 8'b00110110; 
    { 8'hd3, 4'h1 }: pattern = 8'b00110110; 
    { 8'hd3, 4'h2 }: pattern = 8'b00110110; 
    { 8'hd3, 4'h3 }: pattern = 8'b00110110; 
    { 8'hd3, 4'h4 }: pattern = 8'b00110110; 
    { 8'hd3, 4'h5 }: pattern = 8'b00110110; 
    { 8'hd3, 4'h6 }: pattern = 8'b00110110; 
    { 8'hd3, 4'h7 }: pattern = 8'b00111111; 
    { 8'hd3, 4'h8 }: pattern = 8'b00000000; 
    { 8'hd3, 4'h9 }: pattern = 8'b00000000; 
    { 8'hd3, 4'ha }: pattern = 8'b00000000; 
    { 8'hd3, 4'hb }: pattern = 8'b00000000; 
    { 8'hd3, 4'hc }: pattern = 8'b00000000; 
    { 8'hd3, 4'hd }: pattern = 8'b00000000; 
    { 8'hd3, 4'he }: pattern = 8'b00000000; 
    { 8'hd3, 4'hf }: pattern = 8'b00000000; 

    { 8'hd4, 4'h0 }: pattern = 8'b00011000; 
    { 8'hd4, 4'h1 }: pattern = 8'b00011000; 
    { 8'hd4, 4'h2 }: pattern = 8'b00011000; 
    { 8'hd4, 4'h3 }: pattern = 8'b00011000; 
    { 8'hd4, 4'h4 }: pattern = 8'b00011000; 
    { 8'hd4, 4'h5 }: pattern = 8'b00011111; 
    { 8'hd4, 4'h6 }: pattern = 8'b00011000; 
    { 8'hd4, 4'h7 }: pattern = 8'b00011111; 
    { 8'hd4, 4'h8 }: pattern = 8'b00000000; 
    { 8'hd4, 4'h9 }: pattern = 8'b00000000; 
    { 8'hd4, 4'ha }: pattern = 8'b00000000; 
    { 8'hd4, 4'hb }: pattern = 8'b00000000; 
    { 8'hd4, 4'hc }: pattern = 8'b00000000; 
    { 8'hd4, 4'hd }: pattern = 8'b00000000; 
    { 8'hd4, 4'he }: pattern = 8'b00000000; 
    { 8'hd4, 4'hf }: pattern = 8'b00000000; 

    { 8'hd5, 4'h0 }: pattern = 8'b00000000; 
    { 8'hd5, 4'h1 }: pattern = 8'b00000000; 
    { 8'hd5, 4'h2 }: pattern = 8'b00000000; 
    { 8'hd5, 4'h3 }: pattern = 8'b00000000; 
    { 8'hd5, 4'h4 }: pattern = 8'b00000000; 
    { 8'hd5, 4'h5 }: pattern = 8'b00011111; 
    { 8'hd5, 4'h6 }: pattern = 8'b00011000; 
    { 8'hd5, 4'h7 }: pattern = 8'b00011111; 
    { 8'hd5, 4'h8 }: pattern = 8'b00011000; 
    { 8'hd5, 4'h9 }: pattern = 8'b00011000; 
    { 8'hd5, 4'ha }: pattern = 8'b00011000; 
    { 8'hd5, 4'hb }: pattern = 8'b00011000; 
    { 8'hd5, 4'hc }: pattern = 8'b00011000; 
    { 8'hd5, 4'hd }: pattern = 8'b00011000; 
    { 8'hd5, 4'he }: pattern = 8'b00011000; 
    { 8'hd5, 4'hf }: pattern = 8'b00011000; 

    { 8'hd6, 4'h0 }: pattern = 8'b00000000; 
    { 8'hd6, 4'h1 }: pattern = 8'b00000000; 
    { 8'hd6, 4'h2 }: pattern = 8'b00000000; 
    { 8'hd6, 4'h3 }: pattern = 8'b00000000; 
    { 8'hd6, 4'h4 }: pattern = 8'b00000000; 
    { 8'hd6, 4'h5 }: pattern = 8'b00000000; 
    { 8'hd6, 4'h6 }: pattern = 8'b00000000; 
    { 8'hd6, 4'h7 }: pattern = 8'b00111111; 
    { 8'hd6, 4'h8 }: pattern = 8'b00110110; 
    { 8'hd6, 4'h9 }: pattern = 8'b00110110; 
    { 8'hd6, 4'ha }: pattern = 8'b00110110; 
    { 8'hd6, 4'hb }: pattern = 8'b00110110; 
    { 8'hd6, 4'hc }: pattern = 8'b00110110; 
    { 8'hd6, 4'hd }: pattern = 8'b00110110; 
    { 8'hd6, 4'he }: pattern = 8'b00110110; 
    { 8'hd6, 4'hf }: pattern = 8'b00110110; 

    { 8'hd7, 4'h0 }: pattern = 8'b00110110; 
    { 8'hd7, 4'h1 }: pattern = 8'b00110110; 
    { 8'hd7, 4'h2 }: pattern = 8'b00110110; 
    { 8'hd7, 4'h3 }: pattern = 8'b00110110; 
    { 8'hd7, 4'h4 }: pattern = 8'b00110110; 
    { 8'hd7, 4'h5 }: pattern = 8'b00110110; 
    { 8'hd7, 4'h6 }: pattern = 8'b00110110; 
    { 8'hd7, 4'h7 }: pattern = 8'b11111111; 
    { 8'hd7, 4'h8 }: pattern = 8'b00110110; 
    { 8'hd7, 4'h9 }: pattern = 8'b00110110; 
    { 8'hd7, 4'ha }: pattern = 8'b00110110; 
    { 8'hd7, 4'hb }: pattern = 8'b00110110; 
    { 8'hd7, 4'hc }: pattern = 8'b00110110; 
    { 8'hd7, 4'hd }: pattern = 8'b00110110; 
    { 8'hd7, 4'he }: pattern = 8'b00110110; 
    { 8'hd7, 4'hf }: pattern = 8'b00110110; 

    { 8'hd8, 4'h0 }: pattern = 8'b00011000; 
    { 8'hd8, 4'h1 }: pattern = 8'b00011000; 
    { 8'hd8, 4'h2 }: pattern = 8'b00011000; 
    { 8'hd8, 4'h3 }: pattern = 8'b00011000; 
    { 8'hd8, 4'h4 }: pattern = 8'b00011000; 
    { 8'hd8, 4'h5 }: pattern = 8'b11111111; 
    { 8'hd8, 4'h6 }: pattern = 8'b00011000; 
    { 8'hd8, 4'h7 }: pattern = 8'b11111111; 
    { 8'hd8, 4'h8 }: pattern = 8'b00011000; 
    { 8'hd8, 4'h9 }: pattern = 8'b00011000; 
    { 8'hd8, 4'ha }: pattern = 8'b00011000; 
    { 8'hd8, 4'hb }: pattern = 8'b00011000; 
    { 8'hd8, 4'hc }: pattern = 8'b00011000; 
    { 8'hd8, 4'hd }: pattern = 8'b00011000; 
    { 8'hd8, 4'he }: pattern = 8'b00011000; 
    { 8'hd8, 4'hf }: pattern = 8'b00011000; 

    { 8'hd9, 4'h0 }: pattern = 8'b00011000; 
    { 8'hd9, 4'h1 }: pattern = 8'b00011000; 
    { 8'hd9, 4'h2 }: pattern = 8'b00011000; 
    { 8'hd9, 4'h3 }: pattern = 8'b00011000; 
    { 8'hd9, 4'h4 }: pattern = 8'b00011000; 
    { 8'hd9, 4'h5 }: pattern = 8'b00011000; 
    { 8'hd9, 4'h6 }: pattern = 8'b00011000; 
    { 8'hd9, 4'h7 }: pattern = 8'b11111000; 
    { 8'hd9, 4'h8 }: pattern = 8'b00000000; 
    { 8'hd9, 4'h9 }: pattern = 8'b00000000; 
    { 8'hd9, 4'ha }: pattern = 8'b00000000; 
    { 8'hd9, 4'hb }: pattern = 8'b00000000; 
    { 8'hd9, 4'hc }: pattern = 8'b00000000; 
    { 8'hd9, 4'hd }: pattern = 8'b00000000; 
    { 8'hd9, 4'he }: pattern = 8'b00000000; 
    { 8'hd9, 4'hf }: pattern = 8'b00000000; 

    { 8'hda, 4'h0 }: pattern = 8'b00000000; 
    { 8'hda, 4'h1 }: pattern = 8'b00000000; 
    { 8'hda, 4'h2 }: pattern = 8'b00000000; 
    { 8'hda, 4'h3 }: pattern = 8'b00000000; 
    { 8'hda, 4'h4 }: pattern = 8'b00000000; 
    { 8'hda, 4'h5 }: pattern = 8'b00000000; 
    { 8'hda, 4'h6 }: pattern = 8'b00000000; 
    { 8'hda, 4'h7 }: pattern = 8'b00011111; 
    { 8'hda, 4'h8 }: pattern = 8'b00011000; 
    { 8'hda, 4'h9 }: pattern = 8'b00011000; 
    { 8'hda, 4'ha }: pattern = 8'b00011000; 
    { 8'hda, 4'hb }: pattern = 8'b00011000; 
    { 8'hda, 4'hc }: pattern = 8'b00011000; 
    { 8'hda, 4'hd }: pattern = 8'b00011000; 
    { 8'hda, 4'he }: pattern = 8'b00011000; 
    { 8'hda, 4'hf }: pattern = 8'b00011000; 

    { 8'hdb, 4'h0 }: pattern = 8'b11111111; 
    { 8'hdb, 4'h1 }: pattern = 8'b11111111; 
    { 8'hdb, 4'h2 }: pattern = 8'b11111111; 
    { 8'hdb, 4'h3 }: pattern = 8'b11111111; 
    { 8'hdb, 4'h4 }: pattern = 8'b11111111; 
    { 8'hdb, 4'h5 }: pattern = 8'b11111111; 
    { 8'hdb, 4'h6 }: pattern = 8'b11111111; 
    { 8'hdb, 4'h7 }: pattern = 8'b11111111; 
    { 8'hdb, 4'h8 }: pattern = 8'b11111111; 
    { 8'hdb, 4'h9 }: pattern = 8'b11111111; 
    { 8'hdb, 4'ha }: pattern = 8'b11111111; 
    { 8'hdb, 4'hb }: pattern = 8'b11111111; 
    { 8'hdb, 4'hc }: pattern = 8'b11111111; 
    { 8'hdb, 4'hd }: pattern = 8'b11111111; 
    { 8'hdb, 4'he }: pattern = 8'b11111111; 
    { 8'hdb, 4'hf }: pattern = 8'b11111111; 

    { 8'hdc, 4'h0 }: pattern = 8'b00000000; 
    { 8'hdc, 4'h1 }: pattern = 8'b00000000; 
    { 8'hdc, 4'h2 }: pattern = 8'b00000000; 
    { 8'hdc, 4'h3 }: pattern = 8'b00000000; 
    { 8'hdc, 4'h4 }: pattern = 8'b00000000; 
    { 8'hdc, 4'h5 }: pattern = 8'b00000000; 
    { 8'hdc, 4'h6 }: pattern = 8'b00000000; 
    { 8'hdc, 4'h7 }: pattern = 8'b11111111; 
    { 8'hdc, 4'h8 }: pattern = 8'b11111111; 
    { 8'hdc, 4'h9 }: pattern = 8'b11111111; 
    { 8'hdc, 4'ha }: pattern = 8'b11111111; 
    { 8'hdc, 4'hb }: pattern = 8'b11111111; 
    { 8'hdc, 4'hc }: pattern = 8'b11111111; 
    { 8'hdc, 4'hd }: pattern = 8'b11111111; 
    { 8'hdc, 4'he }: pattern = 8'b11111111; 
    { 8'hdc, 4'hf }: pattern = 8'b11111111; 

    { 8'hdd, 4'h0 }: pattern = 8'b11110000; 
    { 8'hdd, 4'h1 }: pattern = 8'b11110000; 
    { 8'hdd, 4'h2 }: pattern = 8'b11110000; 
    { 8'hdd, 4'h3 }: pattern = 8'b11110000; 
    { 8'hdd, 4'h4 }: pattern = 8'b11110000; 
    { 8'hdd, 4'h5 }: pattern = 8'b11110000; 
    { 8'hdd, 4'h6 }: pattern = 8'b11110000; 
    { 8'hdd, 4'h7 }: pattern = 8'b11110000; 
    { 8'hdd, 4'h8 }: pattern = 8'b11110000; 
    { 8'hdd, 4'h9 }: pattern = 8'b11110000; 
    { 8'hdd, 4'ha }: pattern = 8'b11110000; 
    { 8'hdd, 4'hb }: pattern = 8'b11110000; 
    { 8'hdd, 4'hc }: pattern = 8'b11110000; 
    { 8'hdd, 4'hd }: pattern = 8'b11110000; 
    { 8'hdd, 4'he }: pattern = 8'b11110000; 
    { 8'hdd, 4'hf }: pattern = 8'b11110000; 

    { 8'hde, 4'h0 }: pattern = 8'b00001111; 
    { 8'hde, 4'h1 }: pattern = 8'b00001111; 
    { 8'hde, 4'h2 }: pattern = 8'b00001111; 
    { 8'hde, 4'h3 }: pattern = 8'b00001111; 
    { 8'hde, 4'h4 }: pattern = 8'b00001111; 
    { 8'hde, 4'h5 }: pattern = 8'b00001111; 
    { 8'hde, 4'h6 }: pattern = 8'b00001111; 
    { 8'hde, 4'h7 }: pattern = 8'b00001111; 
    { 8'hde, 4'h8 }: pattern = 8'b00001111; 
    { 8'hde, 4'h9 }: pattern = 8'b00001111; 
    { 8'hde, 4'ha }: pattern = 8'b00001111; 
    { 8'hde, 4'hb }: pattern = 8'b00001111; 
    { 8'hde, 4'hc }: pattern = 8'b00001111; 
    { 8'hde, 4'hd }: pattern = 8'b00001111; 
    { 8'hde, 4'he }: pattern = 8'b00001111; 
    { 8'hde, 4'hf }: pattern = 8'b00001111; 

    { 8'hdf, 4'h0 }: pattern = 8'b11111111; 
    { 8'hdf, 4'h1 }: pattern = 8'b11111111; 
    { 8'hdf, 4'h2 }: pattern = 8'b11111111; 
    { 8'hdf, 4'h3 }: pattern = 8'b11111111; 
    { 8'hdf, 4'h4 }: pattern = 8'b11111111; 
    { 8'hdf, 4'h5 }: pattern = 8'b11111111; 
    { 8'hdf, 4'h6 }: pattern = 8'b11111111; 
    { 8'hdf, 4'h7 }: pattern = 8'b00000000; 
    { 8'hdf, 4'h8 }: pattern = 8'b00000000; 
    { 8'hdf, 4'h9 }: pattern = 8'b00000000; 
    { 8'hdf, 4'ha }: pattern = 8'b00000000; 
    { 8'hdf, 4'hb }: pattern = 8'b00000000; 
    { 8'hdf, 4'hc }: pattern = 8'b00000000; 
    { 8'hdf, 4'hd }: pattern = 8'b00000000; 
    { 8'hdf, 4'he }: pattern = 8'b00000000; 
    { 8'hdf, 4'hf }: pattern = 8'b00000000; 

    { 8'he0, 4'h0 }: pattern = 8'b00000000; 
    { 8'he0, 4'h1 }: pattern = 8'b00000000; 
    { 8'he0, 4'h2 }: pattern = 8'b00000000; 
    { 8'he0, 4'h3 }: pattern = 8'b00000000; 
    { 8'he0, 4'h4 }: pattern = 8'b00000000; 
    { 8'he0, 4'h5 }: pattern = 8'b01110110; 
    { 8'he0, 4'h6 }: pattern = 8'b11011100; 
    { 8'he0, 4'h7 }: pattern = 8'b11011000; 
    { 8'he0, 4'h8 }: pattern = 8'b11011000; 
    { 8'he0, 4'h9 }: pattern = 8'b11011000; 
    { 8'he0, 4'ha }: pattern = 8'b11011100; 
    { 8'he0, 4'hb }: pattern = 8'b01110110; 
    { 8'he0, 4'hc }: pattern = 8'b00000000; 
    { 8'he0, 4'hd }: pattern = 8'b00000000; 
    { 8'he0, 4'he }: pattern = 8'b00000000; 
    { 8'he0, 4'hf }: pattern = 8'b00000000; 

    { 8'he1, 4'h0 }: pattern = 8'b00000000; 
    { 8'he1, 4'h1 }: pattern = 8'b00000000; 
    { 8'he1, 4'h2 }: pattern = 8'b01111000; 
    { 8'he1, 4'h3 }: pattern = 8'b11001100; 
    { 8'he1, 4'h4 }: pattern = 8'b11001100; 
    { 8'he1, 4'h5 }: pattern = 8'b11001100; 
    { 8'he1, 4'h6 }: pattern = 8'b11011000; 
    { 8'he1, 4'h7 }: pattern = 8'b11001100; 
    { 8'he1, 4'h8 }: pattern = 8'b11000110; 
    { 8'he1, 4'h9 }: pattern = 8'b11000110; 
    { 8'he1, 4'ha }: pattern = 8'b11000110; 
    { 8'he1, 4'hb }: pattern = 8'b11001100; 
    { 8'he1, 4'hc }: pattern = 8'b00000000; 
    { 8'he1, 4'hd }: pattern = 8'b00000000; 
    { 8'he1, 4'he }: pattern = 8'b00000000; 
    { 8'he1, 4'hf }: pattern = 8'b00000000; 

    { 8'he2, 4'h0 }: pattern = 8'b00000000; 
    { 8'he2, 4'h1 }: pattern = 8'b00000000; 
    { 8'he2, 4'h2 }: pattern = 8'b11111110; 
    { 8'he2, 4'h3 }: pattern = 8'b11000110; 
    { 8'he2, 4'h4 }: pattern = 8'b11000110; 
    { 8'he2, 4'h5 }: pattern = 8'b11000000; 
    { 8'he2, 4'h6 }: pattern = 8'b11000000; 
    { 8'he2, 4'h7 }: pattern = 8'b11000000; 
    { 8'he2, 4'h8 }: pattern = 8'b11000000; 
    { 8'he2, 4'h9 }: pattern = 8'b11000000; 
    { 8'he2, 4'ha }: pattern = 8'b11000000; 
    { 8'he2, 4'hb }: pattern = 8'b11000000; 
    { 8'he2, 4'hc }: pattern = 8'b00000000; 
    { 8'he2, 4'hd }: pattern = 8'b00000000; 
    { 8'he2, 4'he }: pattern = 8'b00000000; 
    { 8'he2, 4'hf }: pattern = 8'b00000000; 

    { 8'he3, 4'h0 }: pattern = 8'b00000000; 
    { 8'he3, 4'h1 }: pattern = 8'b00000000; 
    { 8'he3, 4'h2 }: pattern = 8'b00000000; 
    { 8'he3, 4'h3 }: pattern = 8'b00000000; 
    { 8'he3, 4'h4 }: pattern = 8'b11111110; 
    { 8'he3, 4'h5 }: pattern = 8'b01101100; 
    { 8'he3, 4'h6 }: pattern = 8'b01101100; 
    { 8'he3, 4'h7 }: pattern = 8'b01101100; 
    { 8'he3, 4'h8 }: pattern = 8'b01101100; 
    { 8'he3, 4'h9 }: pattern = 8'b01101100; 
    { 8'he3, 4'ha }: pattern = 8'b01101100; 
    { 8'he3, 4'hb }: pattern = 8'b01101100; 
    { 8'he3, 4'hc }: pattern = 8'b00000000; 
    { 8'he3, 4'hd }: pattern = 8'b00000000; 
    { 8'he3, 4'he }: pattern = 8'b00000000; 
    { 8'he3, 4'hf }: pattern = 8'b00000000; 

    { 8'he4, 4'h0 }: pattern = 8'b00000000; 
    { 8'he4, 4'h1 }: pattern = 8'b00000000; 
    { 8'he4, 4'h2 }: pattern = 8'b00000000; 
    { 8'he4, 4'h3 }: pattern = 8'b11111110; 
    { 8'he4, 4'h4 }: pattern = 8'b11000110; 
    { 8'he4, 4'h5 }: pattern = 8'b01100000; 
    { 8'he4, 4'h6 }: pattern = 8'b00110000; 
    { 8'he4, 4'h7 }: pattern = 8'b00011000; 
    { 8'he4, 4'h8 }: pattern = 8'b00110000; 
    { 8'he4, 4'h9 }: pattern = 8'b01100000; 
    { 8'he4, 4'ha }: pattern = 8'b11000110; 
    { 8'he4, 4'hb }: pattern = 8'b11111110; 
    { 8'he4, 4'hc }: pattern = 8'b00000000; 
    { 8'he4, 4'hd }: pattern = 8'b00000000; 
    { 8'he4, 4'he }: pattern = 8'b00000000; 
    { 8'he4, 4'hf }: pattern = 8'b00000000; 

    { 8'he5, 4'h0 }: pattern = 8'b00000000; 
    { 8'he5, 4'h1 }: pattern = 8'b00000000; 
    { 8'he5, 4'h2 }: pattern = 8'b00000000; 
    { 8'he5, 4'h3 }: pattern = 8'b00000000; 
    { 8'he5, 4'h4 }: pattern = 8'b00000000; 
    { 8'he5, 4'h5 }: pattern = 8'b01111110; 
    { 8'he5, 4'h6 }: pattern = 8'b11011000; 
    { 8'he5, 4'h7 }: pattern = 8'b11011000; 
    { 8'he5, 4'h8 }: pattern = 8'b11011000; 
    { 8'he5, 4'h9 }: pattern = 8'b11011000; 
    { 8'he5, 4'ha }: pattern = 8'b11011000; 
    { 8'he5, 4'hb }: pattern = 8'b01110000; 
    { 8'he5, 4'hc }: pattern = 8'b00000000; 
    { 8'he5, 4'hd }: pattern = 8'b00000000; 
    { 8'he5, 4'he }: pattern = 8'b00000000; 
    { 8'he5, 4'hf }: pattern = 8'b00000000; 

    { 8'he6, 4'h0 }: pattern = 8'b00000000; 
    { 8'he6, 4'h1 }: pattern = 8'b00000000; 
    { 8'he6, 4'h2 }: pattern = 8'b00000000; 
    { 8'he6, 4'h3 }: pattern = 8'b00000000; 
    { 8'he6, 4'h4 }: pattern = 8'b01100110; 
    { 8'he6, 4'h5 }: pattern = 8'b01100110; 
    { 8'he6, 4'h6 }: pattern = 8'b01100110; 
    { 8'he6, 4'h7 }: pattern = 8'b01100110; 
    { 8'he6, 4'h8 }: pattern = 8'b01100110; 
    { 8'he6, 4'h9 }: pattern = 8'b01111100; 
    { 8'he6, 4'ha }: pattern = 8'b01100000; 
    { 8'he6, 4'hb }: pattern = 8'b01100000; 
    { 8'he6, 4'hc }: pattern = 8'b11000000; 
    { 8'he6, 4'hd }: pattern = 8'b00000000; 
    { 8'he6, 4'he }: pattern = 8'b00000000; 
    { 8'he6, 4'hf }: pattern = 8'b00000000; 

    { 8'he7, 4'h0 }: pattern = 8'b00000000; 
    { 8'he7, 4'h1 }: pattern = 8'b00000000; 
    { 8'he7, 4'h2 }: pattern = 8'b00000000; 
    { 8'he7, 4'h3 }: pattern = 8'b00000000; 
    { 8'he7, 4'h4 }: pattern = 8'b01110110; 
    { 8'he7, 4'h5 }: pattern = 8'b11011100; 
    { 8'he7, 4'h6 }: pattern = 8'b00011000; 
    { 8'he7, 4'h7 }: pattern = 8'b00011000; 
    { 8'he7, 4'h8 }: pattern = 8'b00011000; 
    { 8'he7, 4'h9 }: pattern = 8'b00011000; 
    { 8'he7, 4'ha }: pattern = 8'b00011000; 
    { 8'he7, 4'hb }: pattern = 8'b00011000; 
    { 8'he7, 4'hc }: pattern = 8'b00000000; 
    { 8'he7, 4'hd }: pattern = 8'b00000000; 
    { 8'he7, 4'he }: pattern = 8'b00000000; 
    { 8'he7, 4'hf }: pattern = 8'b00000000; 

    { 8'he8, 4'h0 }: pattern = 8'b00000000; 
    { 8'he8, 4'h1 }: pattern = 8'b00000000; 
    { 8'he8, 4'h2 }: pattern = 8'b00000000; 
    { 8'he8, 4'h3 }: pattern = 8'b01111110; 
    { 8'he8, 4'h4 }: pattern = 8'b00011000; 
    { 8'he8, 4'h5 }: pattern = 8'b00111100; 
    { 8'he8, 4'h6 }: pattern = 8'b01100110; 
    { 8'he8, 4'h7 }: pattern = 8'b01100110; 
    { 8'he8, 4'h8 }: pattern = 8'b01100110; 
    { 8'he8, 4'h9 }: pattern = 8'b00111100; 
    { 8'he8, 4'ha }: pattern = 8'b00011000; 
    { 8'he8, 4'hb }: pattern = 8'b01111110; 
    { 8'he8, 4'hc }: pattern = 8'b00000000; 
    { 8'he8, 4'hd }: pattern = 8'b00000000; 
    { 8'he8, 4'he }: pattern = 8'b00000000; 
    { 8'he8, 4'hf }: pattern = 8'b00000000; 

    { 8'he9, 4'h0 }: pattern = 8'b00000000; 
    { 8'he9, 4'h1 }: pattern = 8'b00000000; 
    { 8'he9, 4'h2 }: pattern = 8'b00000000; 
    { 8'he9, 4'h3 }: pattern = 8'b00111000; 
    { 8'he9, 4'h4 }: pattern = 8'b01101100; 
    { 8'he9, 4'h5 }: pattern = 8'b11000110; 
    { 8'he9, 4'h6 }: pattern = 8'b11000110; 
    { 8'he9, 4'h7 }: pattern = 8'b11111110; 
    { 8'he9, 4'h8 }: pattern = 8'b11000110; 
    { 8'he9, 4'h9 }: pattern = 8'b11000110; 
    { 8'he9, 4'ha }: pattern = 8'b01101100; 
    { 8'he9, 4'hb }: pattern = 8'b00111000; 
    { 8'he9, 4'hc }: pattern = 8'b00000000; 
    { 8'he9, 4'hd }: pattern = 8'b00000000; 
    { 8'he9, 4'he }: pattern = 8'b00000000; 
    { 8'he9, 4'hf }: pattern = 8'b00000000; 

    { 8'hea, 4'h0 }: pattern = 8'b00000000; 
    { 8'hea, 4'h1 }: pattern = 8'b00000000; 
    { 8'hea, 4'h2 }: pattern = 8'b00111000; 
    { 8'hea, 4'h3 }: pattern = 8'b01101100; 
    { 8'hea, 4'h4 }: pattern = 8'b11000110; 
    { 8'hea, 4'h5 }: pattern = 8'b11000110; 
    { 8'hea, 4'h6 }: pattern = 8'b11000110; 
    { 8'hea, 4'h7 }: pattern = 8'b01101100; 
    { 8'hea, 4'h8 }: pattern = 8'b01101100; 
    { 8'hea, 4'h9 }: pattern = 8'b01101100; 
    { 8'hea, 4'ha }: pattern = 8'b01101100; 
    { 8'hea, 4'hb }: pattern = 8'b11101110; 
    { 8'hea, 4'hc }: pattern = 8'b00000000; 
    { 8'hea, 4'hd }: pattern = 8'b00000000; 
    { 8'hea, 4'he }: pattern = 8'b00000000; 
    { 8'hea, 4'hf }: pattern = 8'b00000000; 

    { 8'heb, 4'h0 }: pattern = 8'b00000000; 
    { 8'heb, 4'h1 }: pattern = 8'b00000000; 
    { 8'heb, 4'h2 }: pattern = 8'b00011110; 
    { 8'heb, 4'h3 }: pattern = 8'b00110000; 
    { 8'heb, 4'h4 }: pattern = 8'b00011000; 
    { 8'heb, 4'h5 }: pattern = 8'b00001100; 
    { 8'heb, 4'h6 }: pattern = 8'b00111110; 
    { 8'heb, 4'h7 }: pattern = 8'b01100110; 
    { 8'heb, 4'h8 }: pattern = 8'b01100110; 
    { 8'heb, 4'h9 }: pattern = 8'b01100110; 
    { 8'heb, 4'ha }: pattern = 8'b01100110; 
    { 8'heb, 4'hb }: pattern = 8'b00111100; 
    { 8'heb, 4'hc }: pattern = 8'b00000000; 
    { 8'heb, 4'hd }: pattern = 8'b00000000; 
    { 8'heb, 4'he }: pattern = 8'b00000000; 
    { 8'heb, 4'hf }: pattern = 8'b00000000; 

    { 8'hec, 4'h0 }: pattern = 8'b00000000; 
    { 8'hec, 4'h1 }: pattern = 8'b00000000; 
    { 8'hec, 4'h2 }: pattern = 8'b00000000; 
    { 8'hec, 4'h3 }: pattern = 8'b00000000; 
    { 8'hec, 4'h4 }: pattern = 8'b00000000; 
    { 8'hec, 4'h5 }: pattern = 8'b01111110; 
    { 8'hec, 4'h6 }: pattern = 8'b11011011; 
    { 8'hec, 4'h7 }: pattern = 8'b11011011; 
    { 8'hec, 4'h8 }: pattern = 8'b11011011; 
    { 8'hec, 4'h9 }: pattern = 8'b01111110; 
    { 8'hec, 4'ha }: pattern = 8'b00000000; 
    { 8'hec, 4'hb }: pattern = 8'b00000000; 
    { 8'hec, 4'hc }: pattern = 8'b00000000; 
    { 8'hec, 4'hd }: pattern = 8'b00000000; 
    { 8'hec, 4'he }: pattern = 8'b00000000; 
    { 8'hec, 4'hf }: pattern = 8'b00000000; 

    { 8'hed, 4'h0 }: pattern = 8'b00000000; 
    { 8'hed, 4'h1 }: pattern = 8'b00000000; 
    { 8'hed, 4'h2 }: pattern = 8'b00000000; 
    { 8'hed, 4'h3 }: pattern = 8'b00000011; 
    { 8'hed, 4'h4 }: pattern = 8'b00000110; 
    { 8'hed, 4'h5 }: pattern = 8'b01111110; 
    { 8'hed, 4'h6 }: pattern = 8'b11011011; 
    { 8'hed, 4'h7 }: pattern = 8'b11011011; 
    { 8'hed, 4'h8 }: pattern = 8'b11110011; 
    { 8'hed, 4'h9 }: pattern = 8'b01111110; 
    { 8'hed, 4'ha }: pattern = 8'b01100000; 
    { 8'hed, 4'hb }: pattern = 8'b11000000; 
    { 8'hed, 4'hc }: pattern = 8'b00000000; 
    { 8'hed, 4'hd }: pattern = 8'b00000000; 
    { 8'hed, 4'he }: pattern = 8'b00000000; 
    { 8'hed, 4'hf }: pattern = 8'b00000000; 

    { 8'hee, 4'h0 }: pattern = 8'b00000000; 
    { 8'hee, 4'h1 }: pattern = 8'b00000000; 
    { 8'hee, 4'h2 }: pattern = 8'b00011100; 
    { 8'hee, 4'h3 }: pattern = 8'b00110000; 
    { 8'hee, 4'h4 }: pattern = 8'b01100000; 
    { 8'hee, 4'h5 }: pattern = 8'b01100000; 
    { 8'hee, 4'h6 }: pattern = 8'b01111100; 
    { 8'hee, 4'h7 }: pattern = 8'b01100000; 
    { 8'hee, 4'h8 }: pattern = 8'b01100000; 
    { 8'hee, 4'h9 }: pattern = 8'b01100000; 
    { 8'hee, 4'ha }: pattern = 8'b00110000; 
    { 8'hee, 4'hb }: pattern = 8'b00011100; 
    { 8'hee, 4'hc }: pattern = 8'b00000000; 
    { 8'hee, 4'hd }: pattern = 8'b00000000; 
    { 8'hee, 4'he }: pattern = 8'b00000000; 
    { 8'hee, 4'hf }: pattern = 8'b00000000; 

    { 8'hef, 4'h0 }: pattern = 8'b00000000; 
    { 8'hef, 4'h1 }: pattern = 8'b00000000; 
    { 8'hef, 4'h2 }: pattern = 8'b00000000; 
    { 8'hef, 4'h3 }: pattern = 8'b01111100; 
    { 8'hef, 4'h4 }: pattern = 8'b11000110; 
    { 8'hef, 4'h5 }: pattern = 8'b11000110; 
    { 8'hef, 4'h6 }: pattern = 8'b11000110; 
    { 8'hef, 4'h7 }: pattern = 8'b11000110; 
    { 8'hef, 4'h8 }: pattern = 8'b11000110; 
    { 8'hef, 4'h9 }: pattern = 8'b11000110; 
    { 8'hef, 4'ha }: pattern = 8'b11000110; 
    { 8'hef, 4'hb }: pattern = 8'b11000110; 
    { 8'hef, 4'hc }: pattern = 8'b00000000; 
    { 8'hef, 4'hd }: pattern = 8'b00000000; 
    { 8'hef, 4'he }: pattern = 8'b00000000; 
    { 8'hef, 4'hf }: pattern = 8'b00000000; 

    { 8'hf0, 4'h0 }: pattern = 8'b00000000; 
    { 8'hf0, 4'h1 }: pattern = 8'b00000000; 
    { 8'hf0, 4'h2 }: pattern = 8'b00000000; 
    { 8'hf0, 4'h3 }: pattern = 8'b00000000; 
    { 8'hf0, 4'h4 }: pattern = 8'b11111110; 
    { 8'hf0, 4'h5 }: pattern = 8'b00000000; 
    { 8'hf0, 4'h6 }: pattern = 8'b00000000; 
    { 8'hf0, 4'h7 }: pattern = 8'b11111110; 
    { 8'hf0, 4'h8 }: pattern = 8'b00000000; 
    { 8'hf0, 4'h9 }: pattern = 8'b00000000; 
    { 8'hf0, 4'ha }: pattern = 8'b11111110; 
    { 8'hf0, 4'hb }: pattern = 8'b00000000; 
    { 8'hf0, 4'hc }: pattern = 8'b00000000; 
    { 8'hf0, 4'hd }: pattern = 8'b00000000; 
    { 8'hf0, 4'he }: pattern = 8'b00000000; 
    { 8'hf0, 4'hf }: pattern = 8'b00000000; 

    { 8'hf1, 4'h0 }: pattern = 8'b00000000; 
    { 8'hf1, 4'h1 }: pattern = 8'b00000000; 
    { 8'hf1, 4'h2 }: pattern = 8'b00000000; 
    { 8'hf1, 4'h3 }: pattern = 8'b00000000; 
    { 8'hf1, 4'h4 }: pattern = 8'b00011000; 
    { 8'hf1, 4'h5 }: pattern = 8'b00011000; 
    { 8'hf1, 4'h6 }: pattern = 8'b01111110; 
    { 8'hf1, 4'h7 }: pattern = 8'b00011000; 
    { 8'hf1, 4'h8 }: pattern = 8'b00011000; 
    { 8'hf1, 4'h9 }: pattern = 8'b00000000; 
    { 8'hf1, 4'ha }: pattern = 8'b00000000; 
    { 8'hf1, 4'hb }: pattern = 8'b11111111; 
    { 8'hf1, 4'hc }: pattern = 8'b00000000; 
    { 8'hf1, 4'hd }: pattern = 8'b00000000; 
    { 8'hf1, 4'he }: pattern = 8'b00000000; 
    { 8'hf1, 4'hf }: pattern = 8'b00000000; 

    { 8'hf2, 4'h0 }: pattern = 8'b00000000; 
    { 8'hf2, 4'h1 }: pattern = 8'b00000000; 
    { 8'hf2, 4'h2 }: pattern = 8'b00000000; 
    { 8'hf2, 4'h3 }: pattern = 8'b00110000; 
    { 8'hf2, 4'h4 }: pattern = 8'b00011000; 
    { 8'hf2, 4'h5 }: pattern = 8'b00001100; 
    { 8'hf2, 4'h6 }: pattern = 8'b00000110; 
    { 8'hf2, 4'h7 }: pattern = 8'b00001100; 
    { 8'hf2, 4'h8 }: pattern = 8'b00011000; 
    { 8'hf2, 4'h9 }: pattern = 8'b00110000; 
    { 8'hf2, 4'ha }: pattern = 8'b00000000; 
    { 8'hf2, 4'hb }: pattern = 8'b01111110; 
    { 8'hf2, 4'hc }: pattern = 8'b00000000; 
    { 8'hf2, 4'hd }: pattern = 8'b00000000; 
    { 8'hf2, 4'he }: pattern = 8'b00000000; 
    { 8'hf2, 4'hf }: pattern = 8'b00000000; 

    { 8'hf3, 4'h0 }: pattern = 8'b00000000; 
    { 8'hf3, 4'h1 }: pattern = 8'b00000000; 
    { 8'hf3, 4'h2 }: pattern = 8'b00000000; 
    { 8'hf3, 4'h3 }: pattern = 8'b00001100; 
    { 8'hf3, 4'h4 }: pattern = 8'b00011000; 
    { 8'hf3, 4'h5 }: pattern = 8'b00110000; 
    { 8'hf3, 4'h6 }: pattern = 8'b01100000; 
    { 8'hf3, 4'h7 }: pattern = 8'b00110000; 
    { 8'hf3, 4'h8 }: pattern = 8'b00011000; 
    { 8'hf3, 4'h9 }: pattern = 8'b00001100; 
    { 8'hf3, 4'ha }: pattern = 8'b00000000; 
    { 8'hf3, 4'hb }: pattern = 8'b01111110; 
    { 8'hf3, 4'hc }: pattern = 8'b00000000; 
    { 8'hf3, 4'hd }: pattern = 8'b00000000; 
    { 8'hf3, 4'he }: pattern = 8'b00000000; 
    { 8'hf3, 4'hf }: pattern = 8'b00000000; 

    { 8'hf4, 4'h0 }: pattern = 8'b00000000; 
    { 8'hf4, 4'h1 }: pattern = 8'b00000000; 
    { 8'hf4, 4'h2 }: pattern = 8'b00001110; 
    { 8'hf4, 4'h3 }: pattern = 8'b00011011; 
    { 8'hf4, 4'h4 }: pattern = 8'b00011011; 
    { 8'hf4, 4'h5 }: pattern = 8'b00011000; 
    { 8'hf4, 4'h6 }: pattern = 8'b00011000; 
    { 8'hf4, 4'h7 }: pattern = 8'b00011000; 
    { 8'hf4, 4'h8 }: pattern = 8'b00011000; 
    { 8'hf4, 4'h9 }: pattern = 8'b00011000; 
    { 8'hf4, 4'ha }: pattern = 8'b00011000; 
    { 8'hf4, 4'hb }: pattern = 8'b00011000; 
    { 8'hf4, 4'hc }: pattern = 8'b00011000; 
    { 8'hf4, 4'hd }: pattern = 8'b00011000; 
    { 8'hf4, 4'he }: pattern = 8'b00011000; 
    { 8'hf4, 4'hf }: pattern = 8'b00011000; 

    { 8'hf5, 4'h0 }: pattern = 8'b00011000; 
    { 8'hf5, 4'h1 }: pattern = 8'b00011000; 
    { 8'hf5, 4'h2 }: pattern = 8'b00011000; 
    { 8'hf5, 4'h3 }: pattern = 8'b00011000; 
    { 8'hf5, 4'h4 }: pattern = 8'b00011000; 
    { 8'hf5, 4'h5 }: pattern = 8'b00011000; 
    { 8'hf5, 4'h6 }: pattern = 8'b00011000; 
    { 8'hf5, 4'h7 }: pattern = 8'b00011000; 
    { 8'hf5, 4'h8 }: pattern = 8'b11011000; 
    { 8'hf5, 4'h9 }: pattern = 8'b11011000; 
    { 8'hf5, 4'ha }: pattern = 8'b11011000; 
    { 8'hf5, 4'hb }: pattern = 8'b01110000; 
    { 8'hf5, 4'hc }: pattern = 8'b00000000; 
    { 8'hf5, 4'hd }: pattern = 8'b00000000; 
    { 8'hf5, 4'he }: pattern = 8'b00000000; 
    { 8'hf5, 4'hf }: pattern = 8'b00000000; 

    { 8'hf6, 4'h0 }: pattern = 8'b00000000; 
    { 8'hf6, 4'h1 }: pattern = 8'b00000000; 
    { 8'hf6, 4'h2 }: pattern = 8'b00000000; 
    { 8'hf6, 4'h3 }: pattern = 8'b00000000; 
    { 8'hf6, 4'h4 }: pattern = 8'b00011000; 
    { 8'hf6, 4'h5 }: pattern = 8'b00011000; 
    { 8'hf6, 4'h6 }: pattern = 8'b00000000; 
    { 8'hf6, 4'h7 }: pattern = 8'b01111110; 
    { 8'hf6, 4'h8 }: pattern = 8'b00000000; 
    { 8'hf6, 4'h9 }: pattern = 8'b00011000; 
    { 8'hf6, 4'ha }: pattern = 8'b00011000; 
    { 8'hf6, 4'hb }: pattern = 8'b00000000; 
    { 8'hf6, 4'hc }: pattern = 8'b00000000; 
    { 8'hf6, 4'hd }: pattern = 8'b00000000; 
    { 8'hf6, 4'he }: pattern = 8'b00000000; 
    { 8'hf6, 4'hf }: pattern = 8'b00000000; 

    { 8'hf7, 4'h0 }: pattern = 8'b00000000; 
    { 8'hf7, 4'h1 }: pattern = 8'b00000000; 
    { 8'hf7, 4'h2 }: pattern = 8'b00000000; 
    { 8'hf7, 4'h3 }: pattern = 8'b00000000; 
    { 8'hf7, 4'h4 }: pattern = 8'b00000000; 
    { 8'hf7, 4'h5 }: pattern = 8'b01110110; 
    { 8'hf7, 4'h6 }: pattern = 8'b11011100; 
    { 8'hf7, 4'h7 }: pattern = 8'b00000000; 
    { 8'hf7, 4'h8 }: pattern = 8'b01110110; 
    { 8'hf7, 4'h9 }: pattern = 8'b11011100; 
    { 8'hf7, 4'ha }: pattern = 8'b00000000; 
    { 8'hf7, 4'hb }: pattern = 8'b00000000; 
    { 8'hf7, 4'hc }: pattern = 8'b00000000; 
    { 8'hf7, 4'hd }: pattern = 8'b00000000; 
    { 8'hf7, 4'he }: pattern = 8'b00000000; 
    { 8'hf7, 4'hf }: pattern = 8'b00000000; 

    { 8'hf8, 4'h0 }: pattern = 8'b00000000; 
    { 8'hf8, 4'h1 }: pattern = 8'b00111000; 
    { 8'hf8, 4'h2 }: pattern = 8'b01101100; 
    { 8'hf8, 4'h3 }: pattern = 8'b01101100; 
    { 8'hf8, 4'h4 }: pattern = 8'b00111000; 
    { 8'hf8, 4'h5 }: pattern = 8'b00000000; 
    { 8'hf8, 4'h6 }: pattern = 8'b00000000; 
    { 8'hf8, 4'h7 }: pattern = 8'b00000000; 
    { 8'hf8, 4'h8 }: pattern = 8'b00000000; 
    { 8'hf8, 4'h9 }: pattern = 8'b00000000; 
    { 8'hf8, 4'ha }: pattern = 8'b00000000; 
    { 8'hf8, 4'hb }: pattern = 8'b00000000; 
    { 8'hf8, 4'hc }: pattern = 8'b00000000; 
    { 8'hf8, 4'hd }: pattern = 8'b00000000; 
    { 8'hf8, 4'he }: pattern = 8'b00000000; 
    { 8'hf8, 4'hf }: pattern = 8'b00000000; 

    { 8'hf9, 4'h0 }: pattern = 8'b00000000; 
    { 8'hf9, 4'h1 }: pattern = 8'b00000000; 
    { 8'hf9, 4'h2 }: pattern = 8'b00000000; 
    { 8'hf9, 4'h3 }: pattern = 8'b00000000; 
    { 8'hf9, 4'h4 }: pattern = 8'b00000000; 
    { 8'hf9, 4'h5 }: pattern = 8'b00000000; 
    { 8'hf9, 4'h6 }: pattern = 8'b00000000; 
    { 8'hf9, 4'h7 }: pattern = 8'b00011000; 
    { 8'hf9, 4'h8 }: pattern = 8'b00011000; 
    { 8'hf9, 4'h9 }: pattern = 8'b00000000; 
    { 8'hf9, 4'ha }: pattern = 8'b00000000; 
    { 8'hf9, 4'hb }: pattern = 8'b00000000; 
    { 8'hf9, 4'hc }: pattern = 8'b00000000; 
    { 8'hf9, 4'hd }: pattern = 8'b00000000; 
    { 8'hf9, 4'he }: pattern = 8'b00000000; 
    { 8'hf9, 4'hf }: pattern = 8'b00000000; 

    { 8'hfa, 4'h0 }: pattern = 8'b00000000; 
    { 8'hfa, 4'h1 }: pattern = 8'b00000000; 
    { 8'hfa, 4'h2 }: pattern = 8'b00000000; 
    { 8'hfa, 4'h3 }: pattern = 8'b00000000; 
    { 8'hfa, 4'h4 }: pattern = 8'b00000000; 
    { 8'hfa, 4'h5 }: pattern = 8'b00000000; 
    { 8'hfa, 4'h6 }: pattern = 8'b00000000; 
    { 8'hfa, 4'h7 }: pattern = 8'b00000000; 
    { 8'hfa, 4'h8 }: pattern = 8'b00011000; 
    { 8'hfa, 4'h9 }: pattern = 8'b00000000; 
    { 8'hfa, 4'ha }: pattern = 8'b00000000; 
    { 8'hfa, 4'hb }: pattern = 8'b00000000; 
    { 8'hfa, 4'hc }: pattern = 8'b00000000; 
    { 8'hfa, 4'hd }: pattern = 8'b00000000; 
    { 8'hfa, 4'he }: pattern = 8'b00000000; 
    { 8'hfa, 4'hf }: pattern = 8'b00000000; 

    { 8'hfb, 4'h0 }: pattern = 8'b00000000; 
    { 8'hfb, 4'h1 }: pattern = 8'b00001111; 
    { 8'hfb, 4'h2 }: pattern = 8'b00001100; 
    { 8'hfb, 4'h3 }: pattern = 8'b00001100; 
    { 8'hfb, 4'h4 }: pattern = 8'b00001100; 
    { 8'hfb, 4'h5 }: pattern = 8'b00001100; 
    { 8'hfb, 4'h6 }: pattern = 8'b00001100; 
    { 8'hfb, 4'h7 }: pattern = 8'b11101100; 
    { 8'hfb, 4'h8 }: pattern = 8'b01101100; 
    { 8'hfb, 4'h9 }: pattern = 8'b01101100; 
    { 8'hfb, 4'ha }: pattern = 8'b00111100; 
    { 8'hfb, 4'hb }: pattern = 8'b00011100; 
    { 8'hfb, 4'hc }: pattern = 8'b00000000; 
    { 8'hfb, 4'hd }: pattern = 8'b00000000; 
    { 8'hfb, 4'he }: pattern = 8'b00000000; 
    { 8'hfb, 4'hf }: pattern = 8'b00000000; 

    { 8'hfc, 4'h0 }: pattern = 8'b00000000; 
    { 8'hfc, 4'h1 }: pattern = 8'b11011000; 
    { 8'hfc, 4'h2 }: pattern = 8'b01101100; 
    { 8'hfc, 4'h3 }: pattern = 8'b01101100; 
    { 8'hfc, 4'h4 }: pattern = 8'b01101100; 
    { 8'hfc, 4'h5 }: pattern = 8'b01101100; 
    { 8'hfc, 4'h6 }: pattern = 8'b01101100; 
    { 8'hfc, 4'h7 }: pattern = 8'b00000000; 
    { 8'hfc, 4'h8 }: pattern = 8'b00000000; 
    { 8'hfc, 4'h9 }: pattern = 8'b00000000; 
    { 8'hfc, 4'ha }: pattern = 8'b00000000; 
    { 8'hfc, 4'hb }: pattern = 8'b00000000; 
    { 8'hfc, 4'hc }: pattern = 8'b00000000; 
    { 8'hfc, 4'hd }: pattern = 8'b00000000; 
    { 8'hfc, 4'he }: pattern = 8'b00000000; 
    { 8'hfc, 4'hf }: pattern = 8'b00000000; 

    { 8'hfd, 4'h0 }: pattern = 8'b00000000; 
    { 8'hfd, 4'h1 }: pattern = 8'b01110000; 
    { 8'hfd, 4'h2 }: pattern = 8'b11011000; 
    { 8'hfd, 4'h3 }: pattern = 8'b00110000; 
    { 8'hfd, 4'h4 }: pattern = 8'b01100000; 
    { 8'hfd, 4'h5 }: pattern = 8'b11001000; 
    { 8'hfd, 4'h6 }: pattern = 8'b11111000; 
    { 8'hfd, 4'h7 }: pattern = 8'b00000000; 
    { 8'hfd, 4'h8 }: pattern = 8'b00000000; 
    { 8'hfd, 4'h9 }: pattern = 8'b00000000; 
    { 8'hfd, 4'ha }: pattern = 8'b00000000; 
    { 8'hfd, 4'hb }: pattern = 8'b00000000; 
    { 8'hfd, 4'hc }: pattern = 8'b00000000; 
    { 8'hfd, 4'hd }: pattern = 8'b00000000; 
    { 8'hfd, 4'he }: pattern = 8'b00000000; 
    { 8'hfd, 4'hf }: pattern = 8'b00000000; 

    { 8'hfe, 4'h0 }: pattern = 8'b00000000; 
    { 8'hfe, 4'h1 }: pattern = 8'b00000000; 
    { 8'hfe, 4'h2 }: pattern = 8'b00000000; 
    { 8'hfe, 4'h3 }: pattern = 8'b00000000; 
    { 8'hfe, 4'h4 }: pattern = 8'b01111100; 
    { 8'hfe, 4'h5 }: pattern = 8'b01111100; 
    { 8'hfe, 4'h6 }: pattern = 8'b01111100; 
    { 8'hfe, 4'h7 }: pattern = 8'b01111100; 
    { 8'hfe, 4'h8 }: pattern = 8'b01111100; 
    { 8'hfe, 4'h9 }: pattern = 8'b01111100; 
    { 8'hfe, 4'ha }: pattern = 8'b01111100; 
    { 8'hfe, 4'hb }: pattern = 8'b00000000; 
    { 8'hfe, 4'hc }: pattern = 8'b00000000; 
    { 8'hfe, 4'hd }: pattern = 8'b00000000; 
    { 8'hfe, 4'he }: pattern = 8'b00000000; 
    { 8'hfe, 4'hf }: pattern = 8'b00000000; 

    { 8'hff, 4'h0 }: pattern = 8'b00000000; 
    { 8'hff, 4'h1 }: pattern = 8'b00000000; 
    { 8'hff, 4'h2 }: pattern = 8'b00000000; 
    { 8'hff, 4'h3 }: pattern = 8'b00000000; 
    { 8'hff, 4'h4 }: pattern = 8'b00000000; 
    { 8'hff, 4'h5 }: pattern = 8'b00000000; 
    { 8'hff, 4'h6 }: pattern = 8'b00000000; 
    { 8'hff, 4'h7 }: pattern = 8'b00000000; 
    { 8'hff, 4'h8 }: pattern = 8'b00000000; 
    { 8'hff, 4'h9 }: pattern = 8'b00000000; 
    { 8'hff, 4'ha }: pattern = 8'b00000000; 
    { 8'hff, 4'hb }: pattern = 8'b00000000; 
    { 8'hff, 4'hc }: pattern = 8'b00000000; 
    { 8'hff, 4'hd }: pattern = 8'b00000000; 
    { 8'hff, 4'he }: pattern = 8'b00000000; 
    { 8'hff, 4'hf }: pattern = 8'b00000000; 
  endcase

endmodule

